magic
tech sky130A
magscale 1 2
timestamp 1672362834
<< nwell >>
rect 2582 2712 3830 3034
rect 2582 1830 2904 2712
rect 5270 2708 6128 3030
rect 1622 1730 2904 1830
rect 1622 1717 2600 1730
rect 1622 1648 2599 1717
rect 2670 1710 2904 1730
rect 2680 1680 2904 1710
rect 2670 1660 2904 1680
rect 2669 1648 2904 1660
rect 1622 1508 2904 1648
rect 5806 2230 6128 2708
rect 5236 1908 6128 2230
rect 5806 1430 6128 1908
rect 5338 1108 6128 1430
rect 5806 630 6128 1108
rect 5262 620 6128 630
rect 5210 300 6128 620
<< pwell >>
rect 3080 2420 3522 2602
rect 3080 1802 3262 2420
rect 3080 1620 3600 1802
rect 3080 1450 3262 1620
rect 1602 1314 2320 1450
rect 2682 1268 3262 1450
rect 3080 1008 3262 1268
rect 3080 826 3556 1008
rect 3080 216 3262 826
rect 3080 34 3582 216
<< locali >>
rect 3248 2350 3290 2728
rect 3350 2670 3470 2710
rect 3350 2660 3390 2670
rect 5493 2658 5680 2700
rect 5638 2350 5680 2658
rect 3148 2308 5680 2350
rect 2600 1673 2613 1707
rect 2647 1673 2661 1707
rect 2982 1698 3086 1732
rect 3052 1610 3086 1698
rect 3148 1690 3190 2308
rect 3360 2066 3400 2070
rect 3360 2032 3362 2066
rect 3396 2032 3400 2066
rect 3248 1610 3290 1948
rect 3360 1890 3400 2032
rect 3732 1910 3766 1938
rect 3360 1850 3490 1890
rect 5484 1838 5640 1880
rect 2128 1540 2170 1570
rect 3052 1568 3290 1610
rect 2128 1500 2130 1540
rect 3248 1560 3290 1568
rect 5598 1560 5640 1838
rect 3248 1518 5640 1560
rect 2128 1498 2170 1500
rect 2588 1486 2660 1490
rect 2588 1452 2592 1486
rect 2626 1452 2660 1486
rect 2588 1448 2660 1452
rect 2820 1450 3076 1490
rect 3300 1266 3340 1270
rect 3300 1232 3302 1266
rect 3336 1232 3340 1266
rect 3300 1230 3340 1232
rect 3300 1190 3380 1230
rect 3228 990 3270 1128
rect 3340 1090 3380 1190
rect 3340 1050 3500 1090
rect 5486 1038 5660 1080
rect 3230 948 3270 990
rect 3228 760 3270 948
rect 5618 760 5660 1038
rect 3228 718 5660 760
rect 3340 456 3380 460
rect 3340 422 3342 456
rect 3376 422 3380 456
rect 3258 210 3300 318
rect 3340 320 3380 422
rect 3340 280 3490 320
rect 5487 248 5710 290
rect 3170 168 3300 210
rect 3258 -68 3300 168
rect 5668 -68 5710 248
rect 3258 -110 5710 -68
<< viali >>
rect 3248 2728 3290 2770
rect 3732 2738 3766 2772
rect 5180 2660 5230 2710
rect 3350 2620 3390 2660
rect 2613 1673 2647 1707
rect 2948 1698 2982 1732
rect 3362 2032 3396 2066
rect 3148 1648 3190 1690
rect 3248 1948 3290 1990
rect 3732 1938 3766 1972
rect 5180 1850 5230 1900
rect 2130 1500 2170 1540
rect 2242 1462 2276 1496
rect 2592 1452 2626 1486
rect 3076 1450 3110 1490
rect 3302 1232 3336 1266
rect 3228 1128 3270 1170
rect 3722 1138 3756 1172
rect 5180 1060 5230 1110
rect 3188 948 3230 990
rect 3342 422 3376 456
rect 3258 318 3300 360
rect 3722 338 3756 372
rect 3128 168 3170 210
<< metal1 >>
rect 2780 2950 3520 3030
rect 5510 2950 6040 3040
rect 2780 2000 2860 2950
rect 3242 2770 3296 2782
rect 3720 2772 3778 2778
rect 3242 2728 3248 2770
rect 3290 2768 3320 2770
rect 3720 2768 3732 2772
rect 3290 2740 3732 2768
rect 3290 2728 3296 2740
rect 3720 2738 3732 2740
rect 3766 2738 3778 2772
rect 3720 2732 3778 2738
rect 3242 2716 3296 2728
rect 5160 2710 5250 2730
rect 3338 2660 3402 2666
rect 3110 2620 3350 2660
rect 3390 2620 3402 2660
rect 5160 2660 5180 2710
rect 5230 2660 5250 2710
rect 5160 2640 5250 2660
rect 3338 2614 3402 2620
rect 4920 2612 4960 2640
rect 4914 2606 4966 2612
rect 5180 2610 5220 2640
rect 5180 2570 5760 2610
rect 4914 2548 4966 2554
rect 5480 2420 5550 2480
rect 5610 2420 5616 2480
rect 5720 2310 5760 2570
rect 3360 2270 5760 2310
rect 3360 2078 3400 2270
rect 5840 2240 6040 2950
rect 5530 2150 6040 2240
rect 3356 2066 3402 2078
rect 3356 2032 3362 2066
rect 3396 2032 3402 2066
rect 3356 2020 3402 2032
rect 2040 1920 2860 2000
rect 3236 1990 3302 1996
rect 3236 1948 3248 1990
rect 3290 1970 3302 1990
rect 3720 1972 3778 1978
rect 3290 1968 3320 1970
rect 3720 1968 3732 1972
rect 3290 1948 3732 1968
rect 3236 1942 3732 1948
rect 3290 1940 3732 1942
rect 3720 1938 3732 1940
rect 3766 1938 3778 1972
rect 3720 1932 3778 1938
rect 2040 1836 2120 1920
rect 5160 1900 5250 1920
rect 5160 1850 5180 1900
rect 5230 1880 5250 1900
rect 5230 1850 5700 1880
rect 5160 1840 5700 1850
rect 1640 1756 2120 1836
rect 4908 1784 4914 1836
rect 4966 1784 4972 1836
rect 5160 1830 5250 1840
rect 2936 1732 2994 1738
rect 2601 1707 2659 1715
rect 2601 1673 2613 1707
rect 2647 1673 2659 1707
rect 2936 1698 2948 1732
rect 2982 1698 2994 1732
rect 2936 1692 2994 1698
rect 2601 1665 2659 1673
rect 2613 1664 2659 1665
rect 2613 1641 2654 1664
rect 2624 1600 2654 1641
rect 2950 1636 2980 1692
rect 3136 1690 3202 1696
rect 3136 1648 3148 1690
rect 3190 1648 3202 1690
rect 5550 1670 5610 1676
rect 3136 1642 3202 1648
rect 2906 1606 2980 1636
rect 3148 1622 3190 1642
rect 2906 1600 2936 1606
rect 2624 1570 2936 1600
rect 2970 1560 3026 1566
rect 3154 1560 3184 1622
rect 5460 1610 5550 1670
rect 5550 1604 5610 1610
rect 2118 1494 2124 1546
rect 2176 1494 2182 1546
rect 2970 1530 3184 1560
rect 2970 1524 3026 1530
rect 2236 1496 2282 1508
rect 2236 1462 2242 1496
rect 2276 1462 2282 1496
rect 2236 1450 2282 1462
rect 2580 1490 2638 1492
rect 2970 1490 3012 1524
rect 5660 1520 5700 1840
rect 3070 1496 3122 1502
rect 2580 1486 3012 1490
rect 2580 1452 2592 1486
rect 2626 1452 3012 1486
rect 2244 1410 2274 1450
rect 2580 1448 3012 1452
rect 2580 1446 2638 1448
rect 3064 1444 3070 1496
rect 3070 1438 3122 1444
rect 3300 1480 5700 1520
rect 2244 1380 3230 1410
rect 3074 1336 3126 1342
rect 3074 1278 3126 1284
rect 2936 1250 2942 1254
rect 1612 1194 2942 1250
rect 3002 1194 3008 1254
rect 1612 1190 3004 1194
rect 3078 216 3120 1278
rect 3188 1182 3230 1380
rect 3300 1278 3340 1480
rect 5840 1440 6040 2150
rect 5530 1350 6040 1440
rect 3296 1266 3342 1278
rect 3296 1232 3302 1266
rect 3336 1232 3342 1266
rect 3296 1220 3342 1232
rect 3188 1170 3276 1182
rect 3710 1172 3768 1178
rect 3188 1128 3228 1170
rect 3270 1168 3300 1170
rect 3710 1168 3722 1172
rect 3270 1140 3722 1168
rect 3270 1128 3276 1140
rect 3710 1138 3722 1140
rect 3756 1138 3768 1172
rect 3710 1132 3768 1138
rect 3188 1116 3276 1128
rect 3188 1002 3230 1116
rect 5160 1110 5250 1130
rect 5160 1060 5180 1110
rect 5230 1100 5250 1110
rect 5230 1060 5690 1100
rect 5160 1040 5250 1060
rect 3182 990 3236 1002
rect 3182 948 3188 990
rect 3230 948 3236 990
rect 4908 984 4914 1036
rect 4966 984 4972 1036
rect 3182 936 3236 948
rect 5440 810 5550 870
rect 5610 810 5616 870
rect 5650 720 5690 1060
rect 3340 680 5690 720
rect 3340 468 3380 680
rect 5840 640 6040 1350
rect 5540 550 6040 640
rect 3336 456 3382 468
rect 3336 422 3342 456
rect 3376 422 3382 456
rect 3336 410 3382 422
rect 3710 372 3768 378
rect 3252 370 3306 372
rect 3252 368 3330 370
rect 3710 368 3722 372
rect 3252 360 3722 368
rect 3252 318 3258 360
rect 3300 340 3722 360
rect 3300 318 3306 340
rect 3710 338 3722 340
rect 3756 338 3768 372
rect 3710 332 3768 338
rect 3252 306 3306 318
rect 3078 210 3182 216
rect 3078 168 3128 210
rect 3170 168 3182 210
rect 4908 184 4914 236
rect 4966 184 4972 236
rect 3116 162 3182 168
rect 5470 10 5550 70
rect 5610 10 5616 70
rect 5840 10 6040 550
<< via1 >>
rect 4914 2554 4966 2606
rect 5550 2420 5610 2480
rect 4914 1784 4966 1836
rect 5550 1610 5610 1670
rect 2124 1540 2176 1546
rect 2124 1500 2130 1540
rect 2130 1500 2170 1540
rect 2170 1500 2176 1540
rect 2124 1494 2176 1500
rect 3070 1490 3122 1496
rect 3070 1450 3076 1490
rect 3076 1450 3110 1490
rect 3110 1450 3122 1490
rect 3070 1444 3122 1450
rect 3074 1284 3126 1336
rect 2942 1194 3002 1254
rect 4914 984 4966 1036
rect 5550 810 5610 870
rect 4914 184 4966 236
rect 5550 10 5610 70
<< metal2 >>
rect 4908 2554 4914 2606
rect 4966 2554 4972 2606
rect 4920 1842 4960 2554
rect 5560 2486 5700 2490
rect 5550 2480 5700 2486
rect 5610 2420 5700 2480
rect 4914 1836 4966 1842
rect 4914 1778 4966 1784
rect 2124 1546 2176 1552
rect 2124 1488 2176 1494
rect 2128 1410 2170 1488
rect 3064 1444 3070 1496
rect 3122 1490 3128 1496
rect 4920 1490 4960 1778
rect 5550 1670 5700 2420
rect 5544 1610 5550 1670
rect 5610 1610 5700 1670
rect 3122 1450 4960 1490
rect 3122 1444 3128 1450
rect 2128 1368 3010 1410
rect 2970 1330 3010 1368
rect 3068 1330 3074 1336
rect 2970 1290 3074 1330
rect 3068 1284 3074 1290
rect 3126 1284 3132 1336
rect 2942 1254 3002 1260
rect 2942 1186 3002 1194
rect 2942 1126 3080 1186
rect 3020 60 3080 1126
rect 4920 1042 4960 1450
rect 4914 1036 4966 1042
rect 4914 978 4966 984
rect 4920 242 4960 978
rect 5550 870 5700 1610
rect 5610 810 5700 870
rect 4914 236 4966 242
rect 4914 178 4966 184
rect 5550 70 5700 810
rect 3020 10 5550 60
rect 5610 10 5700 70
rect 3020 0 5700 10
use sky130_fd_sc_hd__dfrbp_1  sky130_fd_sc_hd__dfrbp_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1669390400
transform 1 0 3438 0 1 48
box -38 -48 2154 592
use sky130_fd_sc_hd__or4bb_1  sky130_fd_sc_hd__or4bb_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1669390400
transform 1 0 2038 0 1 1248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1669390400
transform 1 0 1604 0 1 1238
box -38 -48 130 592
use sky130_fd_sc_hd__dfrbp_1  x5
timestamp 1669390400
transform 1 0 3438 0 1 2448
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrbp_1  x6
timestamp 1669390400
transform 1 0 3438 0 1 1648
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrbp_1  x7
timestamp 1669390400
transform 1 0 3438 0 1 848
box -38 -48 2154 592
<< labels >>
rlabel locali 5680 -100 5700 -80 1 output
port 2 n
rlabel metal1 3220 2980 3240 3000 1 vcc
port 0 n
rlabel metal1 3150 2630 3170 2650 1 input
port 1 n
rlabel metal2 5620 132 5644 168 1 gnd
port 3 n
<< end >>
