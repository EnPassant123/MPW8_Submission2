magic
tech sky130A
magscale 1 2
timestamp 1671946689
<< pwell >>
rect -201 -5598 201 5598
<< psubdiff >>
rect -165 5528 -69 5562
rect 69 5528 165 5562
rect -165 5466 -131 5528
rect 131 5466 165 5528
rect -165 -5528 -131 -5466
rect 131 -5528 165 -5466
rect -165 -5562 -69 -5528
rect 69 -5562 165 -5528
<< psubdiffcont >>
rect -69 5528 69 5562
rect -165 -5466 -131 5466
rect 131 -5466 165 5466
rect -69 -5562 69 -5528
<< xpolycontact >>
rect -35 5000 35 5432
rect -35 -5432 35 -5000
<< xpolyres >>
rect -35 -5000 35 5000
<< locali >>
rect -165 5528 -69 5562
rect 69 5528 165 5562
rect -165 5466 -131 5528
rect 131 5466 165 5528
rect -165 -5528 -131 -5466
rect 131 -5528 165 -5466
rect -165 -5562 -69 -5528
rect 69 -5562 165 -5528
<< viali >>
rect -19 5017 19 5414
rect -19 -5414 19 -5017
<< metal1 >>
rect -25 5414 25 5426
rect -25 5017 -19 5414
rect 19 5017 25 5414
rect -25 5005 25 5017
rect -25 -5017 25 -5005
rect -25 -5414 -19 -5017
rect 19 -5414 25 -5017
rect -25 -5426 25 -5414
<< res0p35 >>
rect -37 -5002 37 5002
<< properties >>
string FIXED_BBOX -148 -5545 148 5545
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 50 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 286.789k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
