magic
tech sky130A
timestamp 1606063140
<< nwell >>
rect -169 -248 169 248
<< mvpmos >>
rect -40 -100 40 100
<< mvpdiff >>
rect -69 94 -40 100
rect -69 -94 -63 94
rect -46 -94 -40 94
rect -69 -100 -40 -94
rect 40 94 69 100
rect 40 -94 46 94
rect 63 -94 69 94
rect 40 -100 69 -94
<< mvpdiffc >>
rect -63 -94 -46 94
rect 46 -94 63 94
<< mvnsubdiff >>
rect -136 209 136 215
rect -136 192 -82 209
rect 82 192 136 209
rect -136 186 136 192
rect -136 161 -107 186
rect -136 -161 -130 161
rect -113 -161 -107 161
rect 107 161 136 186
rect -136 -186 -107 -161
rect 107 -161 113 161
rect 130 -161 136 161
rect 107 -186 136 -161
rect -136 -192 136 -186
rect -136 -209 -82 -192
rect 82 -209 136 -192
rect -136 -215 136 -209
<< mvnsubdiffcont >>
rect -82 192 82 209
rect -130 -161 -113 161
rect 113 -161 130 161
rect -82 -209 82 -192
<< poly >>
rect -40 140 40 148
rect -40 123 -32 140
rect 32 123 40 140
rect -40 100 40 123
rect -40 -123 40 -100
rect -40 -140 -32 -123
rect 32 -140 40 -123
rect -40 -148 40 -140
<< polycont >>
rect -32 123 32 140
rect -32 -140 32 -123
<< locali >>
rect -130 192 -90 209
rect 90 192 130 209
rect -130 161 -113 192
rect 113 161 130 192
rect -40 123 -32 140
rect 32 123 40 140
rect -63 94 -46 102
rect -63 -102 -46 -94
rect 46 94 63 102
rect 46 -102 63 -94
rect -40 -140 -32 -123
rect 32 -140 40 -123
rect -130 -192 -113 -161
rect 113 -192 130 -161
rect -130 -209 -82 -192
rect 82 -209 130 -192
<< viali >>
rect -90 192 -82 209
rect -82 192 82 209
rect 82 192 90 209
rect -32 123 32 140
rect -63 -94 -46 94
rect 46 -94 63 94
rect -32 -140 32 -123
<< metal1 >>
rect -96 209 96 212
rect -96 192 -90 209
rect 90 192 96 209
rect -96 189 96 192
rect -38 140 38 143
rect -38 123 -32 140
rect 32 123 38 140
rect -38 120 38 123
rect -66 94 -43 100
rect -66 -94 -63 94
rect -46 -94 -43 94
rect -66 -100 -43 -94
rect 43 94 66 100
rect 43 -94 46 94
rect 63 -94 66 94
rect 43 -100 66 -94
rect -38 -123 38 -120
rect -38 -140 -32 -123
rect 32 -140 38 -123
rect -38 -143 38 -140
<< properties >>
string FIXED_BBOX -121 -201 121 201
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 2.00 l 0.80 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 80 viagb 0 viagate 100 viadrn 100 viasrc 100
<< end >>
