magic
tech sky130A
magscale 1 2
timestamp 1672350823
<< pwell >>
rect 313 300 390 550
rect 313 210 390 240
rect 313 200 780 210
rect 313 110 790 200
rect 700 -73 790 110
rect 910 -72 1000 200
<< locali >>
rect -1480 2984 -290 2990
rect -1480 2896 -1474 2984
rect -1386 2896 -290 2984
rect -1480 2890 -290 2896
rect -190 2890 290 2990
rect 390 2890 1310 2990
rect -1270 2770 -1170 2890
rect -870 2880 -830 2890
rect -440 2770 -340 2890
rect 470 2770 570 2890
rect 1190 2780 1290 2890
rect -970 2460 -530 2500
rect -570 2410 -530 2460
rect 620 2430 640 2460
rect 1060 2430 1070 2460
rect -180 2390 270 2430
rect 620 2390 1070 2430
rect 726 2304 815 2310
rect -1360 2030 -1250 2070
rect -785 1955 -715 2225
rect 726 2226 731 2304
rect 809 2226 815 2304
rect 726 2006 815 2226
rect 728 1955 812 2006
rect -785 1885 815 1955
rect -1450 1507 -1410 1510
rect -1450 1473 -1447 1507
rect -1413 1473 -1410 1507
rect -1450 550 -1410 1473
rect -980 680 -940 1780
rect -785 1685 -715 1885
rect -783 1606 -716 1685
rect -783 1537 -716 1539
rect 115 1684 165 1690
rect 115 1646 121 1684
rect 159 1646 165 1684
rect -980 640 -910 680
rect 115 675 165 1646
rect 728 1602 812 1885
rect 970 1740 1070 1780
rect -1450 510 -1180 550
rect -950 390 -910 640
rect -580 630 -140 670
rect -580 390 -540 630
rect 1030 670 1070 1740
rect 380 620 1460 670
rect 745 390 795 620
rect 1560 580 1600 1650
rect 880 577 1600 580
rect 880 543 883 577
rect 917 543 1600 577
rect 880 540 1600 543
rect -960 350 -540 390
rect 570 340 1130 390
rect 230 294 550 300
rect 230 246 496 294
rect 544 246 550 294
rect 230 240 550 246
rect 230 -450 290 240
rect -455 -476 -345 -470
rect -455 -574 -449 -476
rect -351 -574 -345 -476
rect -455 -730 -345 -574
rect 629 -580 670 290
rect -949 -769 -345 -730
rect -800 -770 -345 -769
rect -455 -775 -345 -770
rect 350 -621 670 -580
rect 350 -775 391 -621
rect 629 -670 670 -621
rect -455 -830 425 -775
rect -460 -870 425 -830
rect -455 -885 425 -870
<< viali >>
rect -1474 2896 -1386 2984
rect -290 2890 -190 2990
rect 290 2890 390 2990
rect 1310 2890 1410 2990
rect -785 2225 -715 2295
rect 731 2226 809 2304
rect -1447 1473 -1413 1507
rect -783 1539 -716 1606
rect 121 1646 159 1684
rect 728 1518 812 1602
rect -1180 510 -1140 550
rect 115 625 165 675
rect 1560 1650 1600 1690
rect 883 543 917 577
rect 170 240 230 300
rect 496 246 544 294
rect -449 -574 -351 -476
rect 230 -510 290 -450
rect 425 -885 535 -775
<< metal1 >>
rect -1480 2984 -1380 2996
rect -1480 2896 -1474 2984
rect -1386 2896 -1380 2984
rect -1480 2630 -1380 2896
rect -296 2990 -184 3002
rect -296 2890 -290 2990
rect -190 2890 -184 2990
rect -296 2878 -184 2890
rect 278 2990 402 2996
rect 278 2890 290 2990
rect 390 2890 402 2990
rect 278 2884 402 2890
rect 1304 2990 1416 3002
rect 1304 2890 1310 2990
rect 1410 2890 1416 2990
rect -290 2740 -190 2878
rect -1210 2660 -310 2700
rect -1080 2630 -1040 2660
rect -270 2630 -190 2740
rect -1480 2530 -1210 2630
rect -1310 2210 -1210 2530
rect -1090 2220 -1040 2630
rect -1080 2170 -1040 2220
rect -791 2295 -709 2307
rect -791 2225 -785 2295
rect -715 2290 -709 2295
rect -480 2290 -410 2630
rect -715 2225 -410 2290
rect -791 2220 -410 2225
rect -290 2220 -190 2630
rect 290 2750 390 2884
rect 1304 2878 1416 2890
rect 1310 2750 1410 2878
rect 290 2630 370 2750
rect 400 2660 1300 2720
rect 290 2220 390 2630
rect 500 2310 590 2620
rect 960 2619 1020 2660
rect 1340 2630 1410 2750
rect 1130 2619 1188 2629
rect 960 2560 1190 2619
rect 970 2559 1190 2560
rect 500 2304 821 2310
rect 500 2226 731 2304
rect 809 2226 821 2304
rect 1130 2289 1188 2559
rect 891 2284 1189 2289
rect 500 2220 821 2226
rect 882 2230 1189 2284
rect -791 2213 -709 2220
rect 882 2180 950 2230
rect 1310 2220 1410 2630
rect -1210 2130 -310 2170
rect -1450 1650 -1080 1690
rect -1450 1519 -1410 1650
rect -900 1606 -860 2130
rect 391 2121 1300 2180
rect 109 1684 500 1690
rect -640 1640 -310 1680
rect 109 1646 121 1684
rect 159 1646 500 1684
rect 109 1640 500 1646
rect -795 1610 -704 1612
rect -640 1610 -600 1640
rect -795 1606 -410 1610
rect -1453 1507 -1407 1519
rect -1453 1473 -1447 1507
rect -1413 1473 -1407 1507
rect -1453 1461 -1407 1473
rect -1270 870 -1210 1600
rect -1330 810 -1210 870
rect -1093 1540 -860 1606
rect -1093 1539 -900 1540
rect -800 1539 -783 1606
rect -716 1570 -410 1606
rect -716 1539 -704 1570
rect -1093 817 -1026 1539
rect -795 1533 -704 1539
rect -1330 460 -1270 810
rect -640 770 -600 1570
rect -450 810 -410 1570
rect -290 880 -230 1610
rect 722 1602 818 1614
rect -290 820 -60 880
rect 300 860 390 1600
rect -1180 562 -1140 770
rect -640 730 -310 770
rect -1186 550 -1134 562
rect -1186 510 -1180 550
rect -1140 510 -1134 550
rect -1186 498 -1134 510
rect -120 460 -60 820
rect 0 810 390 860
rect 508 1518 728 1602
rect 812 1518 818 1602
rect 882 1610 941 2121
rect 970 2120 1300 2121
rect 1554 1690 1606 1702
rect 1200 1650 1560 1690
rect 1600 1650 1606 1690
rect 1554 1638 1606 1650
rect 882 1600 1189 1610
rect 882 1551 1190 1600
rect 508 818 592 1518
rect 722 1506 818 1518
rect 1100 820 1190 1551
rect 1300 875 1390 1600
rect 1300 820 1395 875
rect 1305 810 1395 820
rect 0 800 360 810
rect 0 550 60 800
rect 400 760 500 780
rect 120 720 500 760
rect 880 730 1280 770
rect 120 681 160 720
rect 103 675 177 681
rect 103 625 115 675
rect 165 625 177 675
rect 103 619 177 625
rect 880 583 920 730
rect 1340 700 1395 810
rect 871 577 929 583
rect 0 490 390 550
rect 871 543 883 577
rect 917 543 929 577
rect 871 537 929 543
rect 300 465 390 490
rect -1330 400 -60 460
rect 302 453 390 465
rect 1310 453 1395 700
rect -1329 200 -1270 400
rect 302 368 1395 453
rect 164 300 236 312
rect -810 240 170 300
rect 230 240 236 300
rect 164 228 236 240
rect 302 210 390 368
rect 484 294 900 300
rect 484 246 496 294
rect 544 246 900 294
rect 484 240 900 246
rect -860 200 -810 210
rect -1329 141 -810 200
rect -870 -579 -810 141
rect -860 -590 -810 -579
rect -700 -470 -590 210
rect 302 200 780 210
rect 915 200 1025 205
rect 302 112 790 200
rect 218 -450 302 -444
rect -700 -476 -339 -470
rect -700 -574 -449 -476
rect -351 -574 -339 -476
rect 218 -510 230 -450
rect 290 -510 302 -450
rect 218 -516 302 -510
rect -700 -580 -339 -574
rect -700 -590 -650 -580
rect -800 -630 -400 -620
rect 230 -630 290 -516
rect 700 -580 790 112
rect 910 -580 1025 200
rect 915 -600 1025 -580
rect -810 -690 890 -630
rect 940 -720 1025 -600
rect 419 -775 541 -763
rect 915 -775 1025 -720
rect 419 -885 425 -775
rect 535 -885 1025 -775
rect 419 -897 541 -885
use sky130_fd_pr__nfet_01v8_lvt_SMGWK2  XM112
timestamp 1671067782
transform 1 0 446 0 1 1210
box -246 -610 246 610
use sky130_fd_pr__nfet_01v8_lvt_SMGWK2  XM113
timestamp 1671067782
transform 1 0 1246 0 1 1210
box -246 -610 246 610
use sky130_fd_pr__nfet_01v8_lvt_SMGWK2  XM114
timestamp 1671067782
transform 1 0 846 0 1 -190
box -246 -610 246 610
use sky130_fd_pr__nfet_01v8_lvt_SMGWK2  XM117
timestamp 1671067782
transform 1 0 -1154 0 1 1210
box -246 -610 246 610
use sky130_fd_pr__nfet_01v8_lvt_SMGWK2  XM118
timestamp 1671067782
transform 1 0 -354 0 1 1210
box -246 -610 246 610
use sky130_fd_pr__nfet_01v8_lvt_SMGWK2  XM119
timestamp 1671067782
transform 1 0 -754 0 1 -190
box -246 -610 246 610
use sky130_fd_pr__pfet_01v8_lvt_PH9SS5  sky130_fd_pr__pfet_01v8_lvt_PH9SS5_0
timestamp 1672350823
transform 1 0 -1154 0 1 2419
box -246 -419 246 419
use sky130_fd_pr__pfet_01v8_lvt_PH9SS5  sky130_fd_pr__pfet_01v8_lvt_PH9SS5_1
timestamp 1672350823
transform 1 0 -354 0 1 2419
box -246 -419 246 419
use sky130_fd_pr__pfet_01v8_lvt_PH9SS5  sky130_fd_pr__pfet_01v8_lvt_PH9SS5_2
timestamp 1672350823
transform 1 0 446 0 1 2419
box -246 -419 246 419
use sky130_fd_pr__pfet_01v8_lvt_PH9SS5  sky130_fd_pr__pfet_01v8_lvt_PH9SS5_3
timestamp 1672350823
transform 1 0 1246 0 1 2419
box -246 -419 246 419
<< labels >>
rlabel locali -60 -880 0 -820 1 gnd
port 4 n
rlabel locali -1450 1110 -1410 1150 1 voffset
port 2 n
rlabel locali 745 1885 815 1955 1 vout
port 6 n
rlabel locali 1570 1250 1590 1280 1 Vplus
port 1 n
rlabel locali 130 1500 150 1530 1 Vminus
port 3 n
rlabel locali 100 2920 120 2950 1 vdd
port 0 n
rlabel locali 250 10 270 40 1 Nbias
port 5 n
<< end >>
