magic
tech sky130A
timestamp 1671947121
<< nwell >>
rect -123 -609 123 609
<< pmos >>
rect -25 -500 25 500
<< pdiff >>
rect -54 494 -25 500
rect -54 -494 -48 494
rect -31 -494 -25 494
rect -54 -500 -25 -494
rect 25 494 54 500
rect 25 -494 31 494
rect 48 -494 54 494
rect 25 -500 54 -494
<< pdiffc >>
rect -48 -494 -31 494
rect 31 -494 48 494
<< nsubdiff >>
rect -105 574 -57 591
rect 57 574 105 591
rect -105 543 -88 574
rect 88 543 105 574
rect -105 -574 -88 -543
rect 88 -574 105 -543
rect -105 -591 -57 -574
rect 57 -591 105 -574
<< nsubdiffcont >>
rect -57 574 57 591
rect -105 -543 -88 543
rect 88 -543 105 543
rect -57 -591 57 -574
<< poly >>
rect -25 540 25 548
rect -25 523 -17 540
rect 17 523 25 540
rect -25 500 25 523
rect -25 -523 25 -500
rect -25 -540 -17 -523
rect 17 -540 25 -523
rect -25 -548 25 -540
<< polycont >>
rect -17 523 17 540
rect -17 -540 17 -523
<< locali >>
rect -105 574 -57 591
rect 57 574 105 591
rect -105 543 -88 574
rect 88 543 105 574
rect -25 523 -17 540
rect 17 523 25 540
rect -48 494 -31 502
rect -48 -502 -31 -494
rect 31 494 48 502
rect 31 -502 48 -494
rect -25 -540 -17 -523
rect 17 -540 25 -523
rect -105 -574 -88 -543
rect 88 -574 105 -543
rect -105 -591 -57 -574
rect 57 -591 105 -574
<< viali >>
rect -17 523 17 540
rect -48 -494 -31 494
rect 31 -494 48 494
rect -17 -540 17 -523
<< metal1 >>
rect -23 540 23 543
rect -23 523 -17 540
rect 17 523 23 540
rect -23 520 23 523
rect -51 494 -28 500
rect -51 -494 -48 494
rect -31 -494 -28 494
rect -51 -500 -28 -494
rect 28 494 51 500
rect 28 -494 31 494
rect 48 -494 51 494
rect 28 -500 51 -494
rect -23 -523 23 -520
rect -23 -540 -17 -523
rect 17 -540 23 -523
rect -23 -543 23 -540
<< properties >>
string FIXED_BBOX -96 -583 96 583
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 10 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
