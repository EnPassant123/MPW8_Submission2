magic
tech sky130A
magscale 1 2
timestamp 1672362834
<< metal3 >>
rect -13104 12492 -6732 12520
rect -13104 6468 -6816 12492
rect -6752 6468 -6732 12492
rect -13104 6440 -6732 6468
rect -6492 12492 -120 12520
rect -6492 6468 -204 12492
rect -140 6468 -120 12492
rect -6492 6440 -120 6468
rect 120 12492 6492 12520
rect 120 6468 6408 12492
rect 6472 6468 6492 12492
rect 120 6440 6492 6468
rect 6732 12492 13104 12520
rect 6732 6468 13020 12492
rect 13084 6468 13104 12492
rect 6732 6440 13104 6468
rect -13104 6172 -6732 6200
rect -13104 148 -6816 6172
rect -6752 148 -6732 6172
rect -13104 120 -6732 148
rect -6492 6172 -120 6200
rect -6492 148 -204 6172
rect -140 148 -120 6172
rect -6492 120 -120 148
rect 120 6172 6492 6200
rect 120 148 6408 6172
rect 6472 148 6492 6172
rect 120 120 6492 148
rect 6732 6172 13104 6200
rect 6732 148 13020 6172
rect 13084 148 13104 6172
rect 6732 120 13104 148
rect -13104 -148 -6732 -120
rect -13104 -6172 -6816 -148
rect -6752 -6172 -6732 -148
rect -13104 -6200 -6732 -6172
rect -6492 -148 -120 -120
rect -6492 -6172 -204 -148
rect -140 -6172 -120 -148
rect -6492 -6200 -120 -6172
rect 120 -148 6492 -120
rect 120 -6172 6408 -148
rect 6472 -6172 6492 -148
rect 120 -6200 6492 -6172
rect 6732 -148 13104 -120
rect 6732 -6172 13020 -148
rect 13084 -6172 13104 -148
rect 6732 -6200 13104 -6172
rect -13104 -6468 -6732 -6440
rect -13104 -12492 -6816 -6468
rect -6752 -12492 -6732 -6468
rect -13104 -12520 -6732 -12492
rect -6492 -6468 -120 -6440
rect -6492 -12492 -204 -6468
rect -140 -12492 -120 -6468
rect -6492 -12520 -120 -12492
rect 120 -6468 6492 -6440
rect 120 -12492 6408 -6468
rect 6472 -12492 6492 -6468
rect 120 -12520 6492 -12492
rect 6732 -6468 13104 -6440
rect 6732 -12492 13020 -6468
rect 13084 -12492 13104 -6468
rect 6732 -12520 13104 -12492
<< via3 >>
rect -6816 6468 -6752 12492
rect -204 6468 -140 12492
rect 6408 6468 6472 12492
rect 13020 6468 13084 12492
rect -6816 148 -6752 6172
rect -204 148 -140 6172
rect 6408 148 6472 6172
rect 13020 148 13084 6172
rect -6816 -6172 -6752 -148
rect -204 -6172 -140 -148
rect 6408 -6172 6472 -148
rect 13020 -6172 13084 -148
rect -6816 -12492 -6752 -6468
rect -204 -12492 -140 -6468
rect 6408 -12492 6472 -6468
rect 13020 -12492 13084 -6468
<< mimcap >>
rect -13064 12440 -7064 12480
rect -13064 6520 -13024 12440
rect -7104 6520 -7064 12440
rect -13064 6480 -7064 6520
rect -6452 12440 -452 12480
rect -6452 6520 -6412 12440
rect -492 6520 -452 12440
rect -6452 6480 -452 6520
rect 160 12440 6160 12480
rect 160 6520 200 12440
rect 6120 6520 6160 12440
rect 160 6480 6160 6520
rect 6772 12440 12772 12480
rect 6772 6520 6812 12440
rect 12732 6520 12772 12440
rect 6772 6480 12772 6520
rect -13064 6120 -7064 6160
rect -13064 200 -13024 6120
rect -7104 200 -7064 6120
rect -13064 160 -7064 200
rect -6452 6120 -452 6160
rect -6452 200 -6412 6120
rect -492 200 -452 6120
rect -6452 160 -452 200
rect 160 6120 6160 6160
rect 160 200 200 6120
rect 6120 200 6160 6120
rect 160 160 6160 200
rect 6772 6120 12772 6160
rect 6772 200 6812 6120
rect 12732 200 12772 6120
rect 6772 160 12772 200
rect -13064 -200 -7064 -160
rect -13064 -6120 -13024 -200
rect -7104 -6120 -7064 -200
rect -13064 -6160 -7064 -6120
rect -6452 -200 -452 -160
rect -6452 -6120 -6412 -200
rect -492 -6120 -452 -200
rect -6452 -6160 -452 -6120
rect 160 -200 6160 -160
rect 160 -6120 200 -200
rect 6120 -6120 6160 -200
rect 160 -6160 6160 -6120
rect 6772 -200 12772 -160
rect 6772 -6120 6812 -200
rect 12732 -6120 12772 -200
rect 6772 -6160 12772 -6120
rect -13064 -6520 -7064 -6480
rect -13064 -12440 -13024 -6520
rect -7104 -12440 -7064 -6520
rect -13064 -12480 -7064 -12440
rect -6452 -6520 -452 -6480
rect -6452 -12440 -6412 -6520
rect -492 -12440 -452 -6520
rect -6452 -12480 -452 -12440
rect 160 -6520 6160 -6480
rect 160 -12440 200 -6520
rect 6120 -12440 6160 -6520
rect 160 -12480 6160 -12440
rect 6772 -6520 12772 -6480
rect 6772 -12440 6812 -6520
rect 12732 -12440 12772 -6520
rect 6772 -12480 12772 -12440
<< mimcapcontact >>
rect -13024 6520 -7104 12440
rect -6412 6520 -492 12440
rect 200 6520 6120 12440
rect 6812 6520 12732 12440
rect -13024 200 -7104 6120
rect -6412 200 -492 6120
rect 200 200 6120 6120
rect 6812 200 12732 6120
rect -13024 -6120 -7104 -200
rect -6412 -6120 -492 -200
rect 200 -6120 6120 -200
rect 6812 -6120 12732 -200
rect -13024 -12440 -7104 -6520
rect -6412 -12440 -492 -6520
rect 200 -12440 6120 -6520
rect 6812 -12440 12732 -6520
<< metal4 >>
rect -10116 12441 -10012 12640
rect -6836 12492 -6732 12640
rect -13025 12440 -7103 12441
rect -13025 6520 -13024 12440
rect -7104 6520 -7103 12440
rect -13025 6519 -7103 6520
rect -10116 6121 -10012 6519
rect -6836 6468 -6816 12492
rect -6752 6468 -6732 12492
rect -3504 12441 -3400 12640
rect -224 12492 -120 12640
rect -6413 12440 -491 12441
rect -6413 6520 -6412 12440
rect -492 6520 -491 12440
rect -6413 6519 -491 6520
rect -6836 6172 -6732 6468
rect -13025 6120 -7103 6121
rect -13025 200 -13024 6120
rect -7104 200 -7103 6120
rect -13025 199 -7103 200
rect -10116 -199 -10012 199
rect -6836 148 -6816 6172
rect -6752 148 -6732 6172
rect -3504 6121 -3400 6519
rect -224 6468 -204 12492
rect -140 6468 -120 12492
rect 3108 12441 3212 12640
rect 6388 12492 6492 12640
rect 199 12440 6121 12441
rect 199 6520 200 12440
rect 6120 6520 6121 12440
rect 199 6519 6121 6520
rect -224 6172 -120 6468
rect -6413 6120 -491 6121
rect -6413 200 -6412 6120
rect -492 200 -491 6120
rect -6413 199 -491 200
rect -6836 -148 -6732 148
rect -13025 -200 -7103 -199
rect -13025 -6120 -13024 -200
rect -7104 -6120 -7103 -200
rect -13025 -6121 -7103 -6120
rect -10116 -6519 -10012 -6121
rect -6836 -6172 -6816 -148
rect -6752 -6172 -6732 -148
rect -3504 -199 -3400 199
rect -224 148 -204 6172
rect -140 148 -120 6172
rect 3108 6121 3212 6519
rect 6388 6468 6408 12492
rect 6472 6468 6492 12492
rect 9720 12441 9824 12640
rect 13000 12492 13104 12640
rect 6811 12440 12733 12441
rect 6811 6520 6812 12440
rect 12732 6520 12733 12440
rect 6811 6519 12733 6520
rect 6388 6172 6492 6468
rect 199 6120 6121 6121
rect 199 200 200 6120
rect 6120 200 6121 6120
rect 199 199 6121 200
rect -224 -148 -120 148
rect -6413 -200 -491 -199
rect -6413 -6120 -6412 -200
rect -492 -6120 -491 -200
rect -6413 -6121 -491 -6120
rect -6836 -6468 -6732 -6172
rect -13025 -6520 -7103 -6519
rect -13025 -12440 -13024 -6520
rect -7104 -12440 -7103 -6520
rect -13025 -12441 -7103 -12440
rect -10116 -12640 -10012 -12441
rect -6836 -12492 -6816 -6468
rect -6752 -12492 -6732 -6468
rect -3504 -6519 -3400 -6121
rect -224 -6172 -204 -148
rect -140 -6172 -120 -148
rect 3108 -199 3212 199
rect 6388 148 6408 6172
rect 6472 148 6492 6172
rect 9720 6121 9824 6519
rect 13000 6468 13020 12492
rect 13084 6468 13104 12492
rect 13000 6172 13104 6468
rect 6811 6120 12733 6121
rect 6811 200 6812 6120
rect 12732 200 12733 6120
rect 6811 199 12733 200
rect 6388 -148 6492 148
rect 199 -200 6121 -199
rect 199 -6120 200 -200
rect 6120 -6120 6121 -200
rect 199 -6121 6121 -6120
rect -224 -6468 -120 -6172
rect -6413 -6520 -491 -6519
rect -6413 -12440 -6412 -6520
rect -492 -12440 -491 -6520
rect -6413 -12441 -491 -12440
rect -6836 -12640 -6732 -12492
rect -3504 -12640 -3400 -12441
rect -224 -12492 -204 -6468
rect -140 -12492 -120 -6468
rect 3108 -6519 3212 -6121
rect 6388 -6172 6408 -148
rect 6472 -6172 6492 -148
rect 9720 -199 9824 199
rect 13000 148 13020 6172
rect 13084 148 13104 6172
rect 13000 -148 13104 148
rect 6811 -200 12733 -199
rect 6811 -6120 6812 -200
rect 12732 -6120 12733 -200
rect 6811 -6121 12733 -6120
rect 6388 -6468 6492 -6172
rect 199 -6520 6121 -6519
rect 199 -12440 200 -6520
rect 6120 -12440 6121 -6520
rect 199 -12441 6121 -12440
rect -224 -12640 -120 -12492
rect 3108 -12640 3212 -12441
rect 6388 -12492 6408 -6468
rect 6472 -12492 6492 -6468
rect 9720 -6519 9824 -6121
rect 13000 -6172 13020 -148
rect 13084 -6172 13104 -148
rect 13000 -6468 13104 -6172
rect 6811 -6520 12733 -6519
rect 6811 -12440 6812 -6520
rect 12732 -12440 12733 -6520
rect 6811 -12441 12733 -12440
rect 6388 -12640 6492 -12492
rect 9720 -12640 9824 -12441
rect 13000 -12492 13020 -6468
rect 13084 -12492 13104 -6468
rect 13000 -12640 13104 -12492
<< properties >>
string FIXED_BBOX 6732 6440 12812 12520
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 30 l 29.995 val 1.822k carea 2.00 cperi 0.19 nx 4 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
