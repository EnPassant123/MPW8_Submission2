magic
tech sky130A
timestamp 1606502073
<< metal3 >>
rect -1568 1536 1568 1550
rect -1568 -1536 1526 1536
rect 1558 -1536 1568 1536
rect -1568 -1550 1568 -1536
<< via3 >>
rect 1526 -1536 1558 1536
<< mimcap >>
rect -1518 1480 1482 1500
rect -1518 -1480 1166 1480
rect 1462 -1480 1482 1480
rect -1518 -1500 1482 -1480
<< mimcapcontact >>
rect 1166 -1480 1462 1480
<< metal4 >>
rect 1518 1536 1566 1544
rect 1165 1480 1462 1480
rect 1165 -1480 1166 1480
rect 1462 -1480 1462 1480
rect 1165 -1480 1462 -1480
rect 1518 -1536 1526 1536
rect 1558 -1536 1566 1536
rect 1518 -1544 1566 -1536
<< properties >>
string FIXED_BBOX -1568 -1550 1532 1550
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 30.00 l 30.00 val 920.4 carea 1.00 cperi 0.17 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov -10
<< end >>
