magic
tech sky130A
magscale 1 2
timestamp 1672350823
<< error_p >>
rect -34 246 34 247
rect -50 -200 50 -199
<< nwell >>
rect -246 -418 246 418
<< pmoslvt >>
rect -50 -200 50 200
<< pdiff >>
rect -108 188 -50 200
rect -108 -188 -96 188
rect -62 -188 -50 188
rect -108 -200 -50 -188
rect 50 188 108 200
rect 50 -188 62 188
rect 96 -188 108 188
rect 50 -200 108 -188
<< pdiffc >>
rect -96 -188 -62 188
rect 62 -188 96 188
<< nsubdiff >>
rect -210 348 -114 382
rect 114 348 210 382
rect -210 286 -176 348
rect 176 286 210 348
rect -210 -348 -176 -286
rect 176 -348 210 -286
rect -210 -382 -114 -348
rect 114 -382 210 -348
<< nsubdiffcont >>
rect -114 348 114 382
rect -210 -286 -176 286
rect 176 -286 210 286
rect -114 -382 114 -348
<< poly >>
rect -50 280 50 296
rect -50 246 -34 280
rect 34 246 50 280
rect -50 200 50 246
rect -50 -246 50 -200
rect -50 -280 -34 -246
rect 34 -280 50 -246
rect -50 -296 50 -280
<< polycont >>
rect -34 246 34 280
rect -34 -280 34 -246
<< locali >>
rect -210 348 -114 382
rect 114 348 210 382
rect -210 286 -176 348
rect 176 286 210 348
rect -50 246 -34 280
rect 34 246 50 280
rect -96 188 -62 204
rect -96 -204 -62 -188
rect 62 188 96 204
rect 62 -204 96 -188
rect -50 -280 -34 -246
rect 34 -280 50 -246
rect -210 -348 -176 -286
rect 176 -348 210 -286
rect -210 -382 -114 -348
rect 114 -382 210 -348
<< viali >>
rect -34 246 34 280
rect -96 -188 -62 188
rect 62 -188 96 188
rect -34 -280 34 -246
<< metal1 >>
rect -46 280 46 286
rect -46 246 -34 280
rect 34 246 46 280
rect -46 240 46 246
rect -102 188 -56 200
rect -102 -188 -96 188
rect -62 -188 -56 188
rect -102 -200 -56 -188
rect 56 188 102 200
rect 56 -188 62 188
rect 96 -188 102 188
rect 56 -200 102 -188
rect -46 -246 46 -240
rect -46 -280 -34 -246
rect 34 -280 46 -246
rect -46 -286 46 -280
<< properties >>
string FIXED_BBOX -192 -366 192 366
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 2.0 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
