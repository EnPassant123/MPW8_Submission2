magic
tech sky130A
magscale 1 2
timestamp 1672354625
<< error_p >>
rect -29 572 29 578
rect -29 538 -17 572
rect -29 532 29 538
rect -29 -538 29 -532
rect -29 -572 -17 -538
rect -29 -578 29 -572
<< pwell >>
rect -212 -710 212 710
<< nmoslvt >>
rect -16 -500 16 500
<< ndiff >>
rect -74 488 -16 500
rect -74 -488 -62 488
rect -28 -488 -16 488
rect -74 -500 -16 -488
rect 16 488 74 500
rect 16 -488 28 488
rect 62 -488 74 488
rect 16 -500 74 -488
<< ndiffc >>
rect -62 -488 -28 488
rect 28 -488 62 488
<< psubdiff >>
rect -176 640 -80 674
rect 80 640 176 674
rect -176 578 -142 640
rect 142 578 176 640
rect -176 -640 -142 -578
rect 142 -640 176 -578
rect -176 -674 -80 -640
rect 80 -674 176 -640
<< psubdiffcont >>
rect -80 640 80 674
rect -176 -578 -142 578
rect 142 -578 176 578
rect -80 -674 80 -640
<< poly >>
rect -33 572 33 588
rect -33 538 -17 572
rect 17 538 33 572
rect -33 522 33 538
rect -16 500 16 522
rect -16 -522 16 -500
rect -33 -538 33 -522
rect -33 -572 -17 -538
rect 17 -572 33 -538
rect -33 -588 33 -572
<< polycont >>
rect -17 538 17 572
rect -17 -572 17 -538
<< locali >>
rect -176 640 -80 674
rect 80 640 176 674
rect -176 578 -142 640
rect 142 578 176 640
rect -33 538 -17 572
rect 17 538 33 572
rect -62 488 -28 504
rect -62 -504 -28 -488
rect 28 488 62 504
rect 28 -504 62 -488
rect -33 -572 -17 -538
rect 17 -572 33 -538
rect -176 -640 -142 -578
rect 142 -640 176 -578
rect -176 -674 -80 -640
rect 80 -674 176 -640
<< viali >>
rect -17 538 17 572
rect -62 -488 -28 488
rect 28 -488 62 488
rect -17 -572 17 -538
<< metal1 >>
rect -29 572 29 578
rect -29 538 -17 572
rect 17 538 29 572
rect -29 532 29 538
rect -68 488 -22 500
rect -68 -488 -62 488
rect -28 -488 -22 488
rect -68 -500 -22 -488
rect 22 488 68 500
rect 22 -488 28 488
rect 62 -488 68 488
rect 22 -500 68 -488
rect -29 -538 29 -532
rect -29 -572 -17 -538
rect 17 -572 29 -538
rect -29 -578 29 -572
<< properties >>
string FIXED_BBOX -159 -657 159 657
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 5.0 l 0.155 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
