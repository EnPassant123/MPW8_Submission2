magic
tech sky130A
magscale 1 2
timestamp 1672468335
<< metal3 >>
rect -1687 1513 1687 1541
rect -1687 -1513 1603 1513
rect 1667 -1513 1687 1513
rect -1687 -1541 1687 -1513
<< via3 >>
rect 1603 -1513 1667 1513
<< mimcap >>
rect -1647 1461 1355 1501
rect -1647 -1461 -1607 1461
rect 1315 -1461 1355 1461
rect -1647 -1501 1355 -1461
<< mimcapcontact >>
rect -1607 -1461 1315 1461
<< metal4 >>
rect 1587 1513 1683 1529
rect -1608 1461 1316 1462
rect -1608 -1461 -1607 1461
rect 1315 -1461 1316 1461
rect -1608 -1462 1316 -1461
rect 1587 -1513 1603 1513
rect 1667 -1513 1683 1513
rect 1587 -1529 1683 -1513
<< properties >>
string FIXED_BBOX -1687 -1541 1395 1541
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 15.005 l 15.005 val 461.703 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
