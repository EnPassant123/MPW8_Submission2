magic
tech sky130A
magscale 1 2
timestamp 1672477638
<< nwell >>
rect 571575 501082 571896 501689
rect 577196 416028 577701 416358
rect 579552 295479 580051 295800
<< pwell >>
rect 579600 295239 579905 295375
<< locali >>
rect 570957 503354 571553 503355
rect 570957 503321 571514 503354
rect 570957 501035 570991 503321
rect 571517 503205 571553 503320
rect 571517 503175 571551 503205
rect 570957 501001 571559 501035
rect 571025 500945 571273 500951
rect 571025 500899 571031 500945
rect 571077 500899 571273 500945
rect 571025 500893 571273 500899
rect 571525 500849 571559 501001
rect 577280 417704 577402 417758
rect 576760 417657 577402 417704
rect 576580 417651 577402 417657
rect 576580 417540 576586 417651
rect 576697 417596 577402 417651
rect 578354 417633 578959 417703
rect 576697 417578 577374 417596
rect 576697 417540 576971 417578
rect 576580 417534 576971 417540
rect 573874 413492 573996 415916
rect 574670 413498 574792 415922
rect 576329 415889 576371 416322
rect 575472 413464 575594 415888
rect 11832 345340 14054 345380
rect 11832 342944 11872 345340
rect 14014 345172 14054 345340
rect 13980 345166 14318 345172
rect 13980 345118 13986 345166
rect 14034 345118 14318 345166
rect 13980 345112 14318 345118
rect 14014 345096 14054 345112
rect 14083 343567 14133 343701
rect 15499 343589 15617 343809
rect 15499 343483 15505 343589
rect 15611 343483 15617 343589
rect 15499 343477 15617 343483
rect 16221 343201 16416 343311
rect 12442 342530 12556 342630
rect 8430 327681 11417 327795
rect 8430 324773 8544 327681
rect 10827 325073 10941 327681
rect 579723 295745 579889 295779
rect 579544 295430 579790 295470
rect 581399 295365 581667 295539
rect 579723 295201 579887 295235
rect 580943 294997 580977 295235
rect 580913 294963 580977 294997
rect 580913 294127 580947 294963
rect 580913 294093 581003 294127
rect 581930 290484 582210 290490
rect 578460 290070 578500 290300
rect 581930 290216 581936 290484
rect 582204 290216 582210 290484
rect 581930 290070 582210 290216
rect 578460 290030 579470 290070
rect 580050 290030 582210 290070
rect 581930 290008 582210 290030
rect 67688 278647 68501 278748
rect 67688 275741 67789 278647
rect 68400 278457 68501 278647
rect 68400 278368 68405 278457
rect 68496 278368 68501 278457
rect 68400 278362 68501 278368
rect 108725 278415 108895 281131
rect 108725 278245 110589 278415
rect 110759 278245 110760 278415
rect 102515 277437 109119 277443
rect 102515 277399 109075 277437
rect 109113 277399 109119 277437
rect 102515 277393 109119 277399
rect 67688 275640 67844 275741
rect 67743 273428 67844 275640
rect 102515 266667 102565 277393
rect 104482 275836 107864 275916
rect 107784 275569 107864 275836
rect 111993 273311 112043 273317
rect 111993 273273 111999 273311
rect 112037 273273 112043 273311
rect 111620 272574 111720 273156
rect 111620 272486 111626 272574
rect 111714 272486 111720 272574
rect 111620 272480 111720 272486
rect 111993 272485 112043 273273
rect 108629 271578 108679 271599
rect 105745 270569 105795 270575
rect 105745 270531 105751 270569
rect 105789 270531 105795 270569
rect 105745 269791 105795 270531
rect 108584 269590 108754 271578
rect 108424 267274 108924 267308
rect 108424 266786 108430 267274
rect 108918 266786 108924 267274
rect 108424 266780 108924 266786
rect 91371 266617 102565 266667
rect 34446 264092 35292 264196
rect 34446 257118 34550 264092
rect 87000 260446 87441 260504
rect 87499 260446 87538 260504
rect 35514 260107 36830 260113
rect 35514 260025 36743 260107
rect 36824 260025 36830 260107
rect 35514 260020 36830 260025
rect 35514 257348 35607 260020
rect 35713 258553 36239 258555
rect 35713 258519 36203 258553
rect 36237 258519 36239 258553
rect 35713 258517 36239 258519
rect 34446 257026 34452 257118
rect 34544 257026 34550 257118
rect 34446 257020 34550 257026
rect 35847 256244 35893 258517
rect 91371 256693 91421 266617
rect 165684 257239 166336 257339
rect 168014 257239 168828 257339
rect 35847 256210 35853 256244
rect 35887 256210 35893 256244
rect 167755 256234 168887 256304
rect 35847 256204 35893 256210
rect 36328 256142 36548 256146
rect 36220 256042 36548 256142
rect 36220 255966 36324 256042
rect 85619 255997 86553 256083
rect 85619 255985 86461 255997
rect 36220 255874 36226 255966
rect 36318 255874 36324 255966
rect 86455 255911 86461 255985
rect 86547 255911 86553 255997
rect 86455 255905 86553 255911
rect 36220 255868 36324 255874
rect 167309 255503 167433 255553
rect 168828 255244 168870 255284
rect 166813 253568 166923 253651
rect 166813 253470 166819 253568
rect 166917 253470 166923 253568
rect 166813 253464 166923 253470
rect 167343 253340 167453 253574
rect 86327 252773 87295 252855
rect 86327 251393 86409 252773
rect 86129 251311 87375 251393
rect 86129 251303 86409 251311
rect 85639 251269 86409 251303
rect 85639 251229 86331 251269
rect 85639 251221 86255 251229
rect 86249 251159 86255 251221
rect 86325 251159 86331 251229
rect 86249 251153 86331 251159
rect 165684 250844 166128 250944
rect 167777 249826 169205 249896
rect 165564 249032 165874 249072
rect 167237 248931 167449 248981
rect 167237 248053 167287 248931
rect 167137 248003 167287 248053
rect 168844 247516 168884 248526
rect 168844 247476 169596 247516
rect 167185 247040 167295 247147
rect 123055 236789 123279 236847
rect 123055 236674 123113 236789
rect 124203 236723 124419 236781
rect 124203 236674 124261 236723
rect 125257 236691 126497 236749
rect 125257 236674 125315 236691
rect 121075 236616 125315 236674
rect 121075 235955 121133 236616
rect 85756 228275 85802 235679
rect 85295 228229 85802 228275
rect 168339 208129 168681 223073
rect 195296 214992 197744 215334
rect 196223 208129 196565 214992
rect 168339 207787 196565 208129
<< viali >>
rect 571514 503320 571554 503354
rect 571482 501440 571626 501586
rect 571031 500899 571077 500945
rect 571273 500893 571331 500951
rect 571525 500741 571559 500775
rect 576586 417540 576697 417651
rect 578959 417215 579473 417729
rect 576326 415684 576374 415732
rect 13986 345118 14034 345166
rect 13491 343531 13561 343601
rect 14083 343517 14133 343567
rect 15505 343483 15611 343589
rect 16230 343090 16314 343178
rect 11832 342904 11872 342944
rect 2254 337974 2630 338350
rect 10827 324959 10941 325073
rect 579504 295430 579544 295470
rect 581667 295365 581841 295539
rect 581003 294093 581037 294127
rect 578460 290300 578500 290340
rect 581936 290216 582204 290484
rect 68405 278368 68496 278457
rect 110589 278245 110759 278415
rect 109075 277399 109113 277437
rect 70087 268250 70176 268339
rect 83591 268244 83692 268345
rect 104402 275836 104482 275916
rect 111999 273273 112037 273311
rect 111620 273156 111720 273256
rect 111626 272486 111714 272574
rect 111993 272435 112043 272485
rect 105751 270531 105789 270569
rect 105745 269741 105795 269791
rect 108430 266786 108918 267274
rect 87441 260446 87499 260504
rect 36743 260025 36824 260107
rect 35675 258517 35713 258555
rect 36203 258519 36237 258553
rect 34452 257026 34544 257118
rect 91371 256643 91421 256693
rect 35853 256210 35887 256244
rect 168887 256234 168957 256304
rect 36226 255874 36318 255966
rect 86461 255911 86547 255997
rect 167259 255503 167309 255553
rect 166819 253470 166917 253568
rect 81159 251203 81269 251313
rect 86255 251159 86325 251229
rect 169205 249826 169275 249896
rect 165524 249032 165564 249072
rect 167087 248003 167137 248053
rect 169596 247476 169636 247516
rect 87470 241688 87834 242052
rect 121075 235897 121133 235955
rect 89316 235359 89634 235677
rect 85249 228229 85295 228275
rect 168339 223073 168681 223415
<< metal1 >>
rect 571502 503314 571508 503366
rect 571560 503314 571566 503366
rect 571508 503308 571560 503314
rect 571456 501588 571656 501614
rect 572150 501606 572342 501612
rect 571025 501469 571324 501527
rect 571025 500951 571083 501469
rect 571456 501438 571482 501588
rect 571630 501438 571656 501588
rect 571456 501414 571656 501438
rect 571840 501294 571900 501446
rect 572144 501414 572150 501606
rect 572342 501414 572348 501606
rect 572150 501408 572342 501414
rect 571267 500951 571337 500963
rect 571019 500945 571089 500951
rect 571019 500899 571031 500945
rect 571077 500899 571089 500945
rect 571019 500893 571089 500899
rect 571267 500893 571273 500951
rect 571331 500893 571337 500951
rect 571267 500881 571337 500893
rect 571273 500833 571331 500881
rect 571516 500784 571568 500790
rect 571513 500735 571516 500781
rect 571568 500735 571571 500781
rect 571516 500726 571568 500732
rect 568897 497307 568903 497457
rect 569053 497307 569802 497457
rect 573609 496151 573821 496254
rect 573718 496070 573821 496151
rect 573718 495973 576654 496070
rect 573720 495826 576654 495973
rect 576898 495826 576904 496070
rect 568994 494830 569352 494890
rect 568994 494042 569054 494830
rect 582222 494206 582282 494212
rect 582222 494042 582282 494146
rect 568994 493982 582282 494042
rect 577586 449278 582142 449981
rect 582845 449278 582851 449981
rect 15176 430948 15182 431528
rect 15762 430948 15768 431528
rect 15182 425218 15762 430948
rect 24684 430264 24690 431324
rect 25750 430264 25756 431324
rect 20356 427598 20362 428058
rect 20822 427598 20828 428058
rect 20362 427092 20822 427598
rect 24690 426858 25750 430264
rect 577586 427002 578289 449278
rect 22032 425798 25750 426858
rect 15182 424638 17732 425218
rect 576266 424294 576272 424394
rect 576372 424294 577489 424394
rect 578533 422439 578922 422614
rect 579097 422439 579103 422614
rect 576630 417876 576742 417882
rect 576742 417764 577160 417876
rect 576630 417758 576742 417764
rect 578953 417735 579479 417741
rect 576580 417657 576703 417663
rect 576574 417534 576580 417657
rect 576703 417534 576709 417657
rect 576580 417528 576703 417534
rect 578947 417209 578953 417735
rect 579479 417209 579485 417735
rect 578953 417203 579479 417209
rect 27813 417021 28663 417027
rect 22561 416171 27813 417021
rect 27813 416165 28663 416171
rect 572822 416270 573022 416276
rect 576063 416270 576573 416400
rect 573022 416070 573506 416270
rect 576063 416202 577512 416270
rect 576310 416070 577512 416202
rect 572822 416064 573022 416070
rect 576324 416034 576376 416040
rect 576324 415976 576376 415982
rect 576326 415738 576374 415976
rect 576314 415732 576386 415738
rect 576314 415684 576326 415732
rect 576374 415684 576386 415732
rect 576314 415678 576386 415684
rect 576326 415174 576374 415678
rect 576318 415122 576324 415174
rect 576376 415122 576382 415174
rect 578077 415077 578135 415433
rect 576164 415019 578135 415077
rect 576324 414932 576376 414938
rect 576324 414874 576376 414880
rect 15800 414541 17732 414562
rect 15800 413982 15937 414541
rect 16591 413982 17732 414541
rect 15937 413881 16591 413887
rect 576326 413528 576374 414874
rect 575900 413480 576374 413528
rect 573594 413392 573646 413398
rect 573594 413334 573646 413340
rect 573597 413331 573643 413334
rect 576043 413309 576091 413480
rect 19894 413033 20016 413040
rect 19891 412983 20372 413033
rect 19894 412974 20016 412983
rect 19894 412846 20016 412852
rect 20302 410971 20512 411408
rect 20296 410761 20302 410971
rect 20512 410761 20518 410971
rect 9298 371169 9304 371411
rect 9546 371169 9552 371411
rect 9304 369670 9546 371169
rect 9262 340066 9494 363732
rect 22866 362111 225797 363729
rect 13980 345172 14040 345178
rect 13974 345112 13980 345172
rect 14040 345112 14046 345172
rect 13980 345106 14040 345112
rect 11826 342950 11878 342956
rect 11820 342898 11826 342950
rect 11878 342898 11884 342950
rect 11826 342892 11878 342898
rect 12434 342762 12558 345028
rect 13485 343607 13567 343613
rect 13479 343537 13485 343607
rect 13567 343537 13573 343607
rect 15499 343595 15617 343601
rect 13479 343531 13491 343537
rect 13561 343531 13573 343537
rect 13479 343525 13573 343531
rect 14077 343573 14139 343579
rect 14077 343567 14087 343573
rect 14077 343517 14083 343567
rect 14077 343511 14087 343517
rect 14139 343511 14145 343573
rect 14077 343505 14139 343511
rect 15499 343471 15617 343477
rect 16200 343487 16350 344088
rect 18117 343601 18247 343607
rect 16200 343337 16905 343487
rect 18111 343471 18117 343601
rect 18235 343471 18247 343601
rect 18117 343465 18247 343471
rect 16200 343178 16350 343337
rect 16200 343090 16230 343178
rect 16314 343090 16350 343178
rect 16200 343064 16350 343090
rect 9262 339828 9494 339834
rect 10738 342182 12558 342762
rect 16755 342533 16905 343337
rect 2248 338356 2636 338362
rect 2242 337980 2248 338356
rect 2636 337980 2642 338356
rect 2242 337974 2254 337980
rect 2630 337974 2642 337980
rect 2242 337968 2642 337974
rect 10738 337406 11318 342182
rect 12434 342002 12558 342182
rect 13756 341352 13796 342146
rect 16397 341473 17247 342533
rect 14314 341358 14366 341364
rect 13756 341312 14314 341352
rect 14314 341300 14366 341306
rect 16391 340623 16397 341473
rect 17247 340623 17253 341473
rect 10738 333562 14740 337406
rect 18584 333562 18590 337406
rect 10738 329052 11318 333562
rect 22866 332383 24484 362111
rect 22860 330765 22866 332383
rect 24484 330765 24490 332383
rect 12105 330691 12239 330703
rect 12105 330581 12111 330691
rect 12233 330581 12239 330691
rect 123136 330645 129751 330759
rect 129865 330645 129871 330759
rect 12111 330575 12233 330581
rect 4892 328472 11318 329052
rect 4892 322458 5472 328472
rect 12238 328276 12244 328544
rect 12512 328276 12518 328544
rect 12244 328072 12512 328276
rect 7492 327892 7544 327898
rect 8252 327891 9143 328019
rect 7544 327841 9143 327891
rect 7492 327834 7544 327840
rect 8252 327801 9143 327841
rect 10858 327804 12526 328072
rect 8252 327036 8470 327801
rect 10815 325073 10953 325079
rect 10815 324959 10827 325073
rect 10941 324959 10953 325073
rect 10815 324953 10953 324959
rect 10827 324838 10941 324953
rect 11773 324838 12623 324844
rect 6122 323962 6128 324422
rect 6588 323962 8562 324422
rect 9982 323988 11773 324838
rect 11773 323982 12623 323988
rect 8330 311186 8336 311290
rect 8440 311186 8446 311290
rect 8336 310907 8440 311186
rect 8062 310857 8440 310907
rect 8062 310717 8112 310857
rect 8336 310830 8440 310857
rect 7492 308846 7544 308852
rect 8062 308845 8112 309158
rect 7544 308795 8112 308845
rect 7492 308788 7544 308794
rect 10832 308572 11908 308772
rect 4892 308208 5482 308214
rect 4892 307612 5482 307618
rect 11708 306480 11908 308572
rect 11702 306280 11708 306480
rect 11908 306280 11914 306480
rect 102969 289071 104089 289285
rect 102969 288984 104135 289071
rect 102969 288906 104134 288984
rect 102969 288824 104089 288906
rect 111576 288824 111856 288920
rect 102969 288763 104041 288824
rect 113128 288820 113634 288920
rect 113734 288820 113740 288920
rect 102969 285987 103491 288763
rect 107379 287898 107873 288335
rect 111687 288280 111856 288338
rect 113168 288280 113448 288380
rect 113548 288280 113554 288380
rect 107379 287404 109620 287898
rect 109984 287510 109990 287562
rect 110042 287561 110048 287562
rect 110042 287511 110775 287561
rect 110042 287510 110048 287511
rect 109126 286792 109620 287404
rect 109126 286298 109626 286792
rect 102969 285465 108273 285987
rect 109120 285798 109126 286298
rect 109626 285798 109632 286298
rect 35038 276629 35044 276767
rect 35182 276629 35188 276767
rect 35044 270701 35182 276629
rect 67798 276621 67904 278496
rect 68014 278463 68112 278500
rect 68793 278463 68894 278469
rect 68011 278457 68793 278463
rect 68011 278368 68405 278457
rect 68496 278368 68793 278457
rect 68011 278362 68793 278368
rect 68894 278362 70182 278463
rect 67455 276515 67904 276621
rect 68014 276518 68112 278362
rect 68793 278356 68894 278362
rect 67455 276055 67561 276515
rect 67798 276512 67904 276515
rect 69939 276458 69993 276464
rect 67882 276404 69939 276458
rect 69993 276404 70002 276458
rect 69939 276398 69993 276404
rect 67449 275949 67455 276055
rect 67561 275949 67567 276055
rect 67455 275621 67561 275949
rect 70081 275779 70182 278362
rect 70495 276458 70549 276464
rect 70362 276404 70495 276458
rect 70549 276404 70927 276458
rect 70495 276398 70549 276404
rect 67455 275515 67927 275621
rect 67821 273637 67927 275515
rect 68044 273755 68152 275628
rect 68547 273755 68657 273761
rect 68042 273645 68547 273755
rect 68044 273636 68152 273645
rect 68261 273639 68657 273645
rect 67892 273528 68050 273580
rect 66047 273405 66849 273411
rect 66849 273320 67505 273405
rect 67892 273320 67944 273528
rect 66849 273268 67944 273320
rect 66849 272603 67505 273268
rect 66047 272597 66849 272603
rect 68261 267691 68591 273639
rect 69825 268603 70439 275779
rect 70873 272773 70927 276404
rect 102969 275999 103491 285465
rect 108180 284929 108230 285465
rect 108894 284224 108900 284276
rect 108952 284224 108958 284276
rect 108901 284095 108951 284224
rect 107588 283926 107640 283932
rect 107588 283868 107640 283874
rect 109464 283814 109470 283866
rect 109522 283814 109528 283866
rect 110725 282530 110775 287511
rect 111114 287550 111166 287556
rect 111166 287499 112959 287549
rect 111114 287492 111166 287498
rect 108227 282156 108277 282530
rect 110223 282480 110775 282530
rect 108220 282104 108226 282156
rect 108278 282104 108284 282156
rect 108471 280076 108521 280960
rect 108470 280070 108522 280076
rect 108470 280012 108522 280018
rect 102969 275869 102999 275999
rect 103129 275916 103491 275999
rect 104884 279839 106750 279980
rect 104396 275916 104488 275928
rect 103129 275869 104402 275916
rect 102969 275836 104402 275869
rect 104482 275836 104488 275916
rect 69819 267989 69825 268603
rect 70439 267989 70445 268603
rect 68255 267361 68261 267691
rect 68591 267361 68597 267691
rect 70870 267294 70931 272773
rect 87108 268636 87244 268642
rect 83328 267989 83334 268603
rect 83948 267989 83954 268603
rect 70836 267288 70968 267294
rect 70968 267156 70970 267288
rect 70836 267150 70968 267156
rect 36691 264895 36697 264988
rect 36790 264895 36796 264988
rect 35056 263577 35149 264738
rect 36697 263577 36790 264895
rect 35056 263484 79440 263577
rect 36747 260380 36840 260388
rect 34962 260258 36064 260342
rect 34962 259944 35046 260258
rect 35297 260017 35683 260087
rect 34962 259860 35272 259944
rect 35188 258968 35272 259860
rect 35392 259847 35462 259950
rect 35613 259847 35683 260017
rect 35392 259777 35683 259847
rect 35392 259063 35462 259777
rect 35392 258993 35731 259063
rect 35392 258970 35462 258993
rect 35661 258909 35731 258993
rect 35980 258972 36064 260258
rect 36737 260287 37439 260380
rect 37532 260287 37538 260380
rect 36737 260113 36830 260287
rect 36731 260107 36836 260113
rect 36731 260025 36743 260107
rect 36824 260025 36836 260107
rect 36731 260019 36836 260025
rect 36210 258972 36294 259872
rect 36416 259870 36508 259872
rect 36737 259870 36830 260019
rect 36415 259777 36830 259870
rect 33477 258839 33483 258909
rect 33553 258839 35731 258909
rect 35558 258758 35564 258764
rect 35254 258718 35564 258758
rect 35254 258616 35294 258718
rect 35558 258712 35564 258718
rect 35616 258712 35622 258764
rect 35252 258576 35414 258616
rect 35661 258555 35731 258839
rect 35964 258888 36294 258972
rect 35778 258764 35830 258770
rect 35964 258758 36048 258888
rect 36416 258884 36508 259777
rect 36926 258900 37050 258902
rect 36926 258840 49864 258900
rect 36312 258794 49864 258840
rect 35830 258718 36048 258758
rect 36926 258744 49864 258794
rect 50020 258744 50026 258900
rect 36926 258742 37050 258744
rect 35778 258706 35830 258712
rect 35964 258708 36048 258718
rect 35174 257624 35278 258530
rect 35661 258522 35675 258555
rect 35014 257520 35278 257624
rect 35388 258517 35675 258522
rect 35713 258517 35731 258555
rect 35388 258452 35731 258517
rect 35964 258624 36754 258708
rect 35388 257542 35458 258452
rect 35964 258280 36048 258624
rect 36191 258553 36249 258559
rect 36191 258519 36203 258553
rect 36237 258519 36249 258553
rect 36191 258513 36249 258519
rect 36670 258518 36754 258624
rect 37508 258518 37592 258524
rect 36201 258360 36239 258513
rect 36670 258434 37508 258518
rect 37508 258428 37592 258434
rect 36201 258322 36436 258360
rect 35964 258196 36302 258280
rect 34446 257124 34550 257130
rect 35014 257124 35118 257520
rect 34446 257118 35118 257124
rect 34446 257026 34452 257118
rect 34544 257026 35118 257118
rect 34446 257020 35118 257026
rect 34446 257014 34550 257020
rect 35014 255972 35118 257020
rect 36218 256298 36302 258196
rect 36420 256402 36522 258278
rect 36418 256298 36778 256402
rect 35847 256250 35893 256256
rect 35847 256244 36462 256250
rect 35847 256210 35853 256244
rect 35887 256210 36462 256244
rect 35847 256204 36462 256210
rect 35847 256198 35893 256204
rect 36220 255972 36324 255978
rect 36674 255972 36778 256298
rect 37218 255972 37322 255974
rect 35014 255966 37354 255972
rect 35014 255874 36226 255966
rect 36318 255874 37354 255966
rect 35014 255868 37354 255874
rect 35448 255778 36082 255868
rect 36220 255862 36324 255868
rect 37218 255282 37322 255868
rect 38630 255282 38734 255288
rect 37218 255178 38630 255282
rect 38630 255172 38734 255178
rect 35448 255138 36082 255144
rect 79347 235311 79440 263484
rect 83334 258830 83948 267989
rect 87108 267006 87244 268500
rect 102969 267629 103491 275836
rect 104396 275824 104488 275836
rect 104884 270470 105025 279839
rect 108620 276371 108670 279930
rect 109660 279880 112043 279930
rect 111330 279072 111382 279078
rect 109069 279021 111330 279071
rect 109069 277727 109119 279021
rect 111330 279014 111382 279020
rect 110583 278421 110765 278427
rect 110583 278415 110595 278421
rect 110583 278245 110589 278415
rect 110583 278239 110595 278245
rect 110765 278239 110771 278421
rect 110583 278233 110765 278239
rect 108979 277489 109153 277727
rect 108973 277315 108979 277489
rect 109153 277315 109159 277489
rect 105745 276321 108670 276371
rect 105745 270569 105795 276321
rect 109069 276114 109119 277315
rect 109068 276014 111720 276114
rect 107805 275869 107811 275999
rect 107941 275869 107947 275999
rect 107811 275494 107941 275869
rect 108534 275830 108586 275836
rect 109069 275829 109119 276014
rect 108586 275779 109119 275829
rect 108534 275772 108586 275778
rect 107253 275364 109125 275494
rect 108534 275098 108586 275104
rect 108534 275040 108586 275046
rect 108535 274534 108585 275040
rect 107556 274328 107562 274380
rect 107614 274328 107620 274380
rect 109460 274268 109466 274320
rect 109518 274268 109524 274320
rect 111620 273262 111720 276014
rect 111993 273311 112043 279880
rect 111993 273273 111999 273311
rect 112037 273273 112043 273311
rect 111608 273256 111732 273262
rect 111993 273261 112043 273273
rect 111608 273156 111620 273256
rect 111720 273156 111732 273256
rect 111608 273150 111732 273156
rect 108080 272985 108132 272991
rect 112909 272984 112959 287499
rect 114920 287348 115400 287354
rect 114914 286880 114920 287348
rect 115400 286880 115406 287348
rect 114914 286868 115406 286880
rect 110181 272934 112959 272984
rect 108080 272927 108132 272933
rect 111620 272580 111720 272586
rect 111614 272480 111620 272580
rect 111720 272480 111726 272580
rect 111981 272485 112055 272491
rect 111620 272474 111720 272480
rect 111981 272435 111993 272485
rect 112043 272435 112055 272485
rect 111981 272429 112055 272435
rect 108425 271122 108475 271414
rect 108418 271070 108424 271122
rect 108476 271070 108482 271122
rect 105745 270531 105751 270569
rect 105789 270531 105795 270569
rect 105745 270519 105795 270531
rect 104884 270329 106752 270470
rect 104884 269400 105035 270329
rect 105739 269791 105801 269803
rect 108543 269791 108593 270405
rect 111993 270377 112043 272429
rect 109597 270327 112043 270377
rect 105739 269741 105745 269791
rect 105795 269741 108593 269791
rect 105739 269729 105801 269741
rect 104878 269296 104884 269400
rect 104988 269296 105035 269400
rect 104894 269290 105035 269296
rect 91419 267107 103491 267629
rect 91419 267086 103381 267107
rect 88653 260959 88983 260965
rect 87963 260931 88653 260959
rect 87061 260629 88653 260931
rect 88983 260629 89300 260931
rect 87061 260601 89300 260629
rect 87435 260510 87505 260516
rect 87435 260504 87447 260510
rect 87435 260446 87441 260504
rect 87435 260440 87447 260446
rect 87505 260440 87511 260510
rect 87435 260434 87505 260440
rect 82416 258160 87130 258830
rect 91419 258160 91945 267086
rect 107009 266519 107059 269741
rect 108424 267280 108924 267286
rect 108418 266780 108424 267280
rect 108924 266780 108930 267280
rect 108424 266774 108924 266780
rect 82416 257638 91945 258160
rect 92529 266469 107059 266519
rect 82416 257530 87130 257638
rect 81147 251313 81281 251319
rect 81147 251307 81159 251313
rect 81269 251307 81281 251313
rect 81147 251197 81153 251307
rect 81275 251197 81281 251307
rect 81153 251191 81275 251197
rect 79968 239428 81268 239434
rect 82416 239428 83716 257530
rect 86505 256003 86603 257530
rect 91359 256637 91365 256699
rect 91417 256693 91433 256699
rect 91421 256643 91433 256693
rect 91417 256637 91433 256643
rect 86211 255997 87207 256003
rect 85675 255884 85898 255918
rect 86211 255911 86461 255997
rect 86547 255911 87207 255997
rect 86211 255905 87207 255911
rect 85675 255826 85709 255884
rect 86211 255828 86309 255905
rect 85675 255770 85744 255826
rect 85675 255250 85742 255770
rect 85870 255730 86309 255828
rect 85675 255189 85709 255250
rect 85870 255246 85968 255730
rect 87109 255455 87207 255905
rect 90578 255694 90584 256002
rect 90892 255694 90898 256002
rect 85675 255155 85843 255189
rect 85675 254797 85709 255155
rect 85339 254623 85345 254797
rect 85519 254623 85836 254797
rect 85662 253922 85836 254623
rect 87093 252715 87211 253363
rect 86811 252597 87211 252715
rect 86811 252561 86929 252597
rect 90584 252561 90892 255694
rect 92529 253213 92579 266469
rect 91225 253163 92579 253213
rect 91225 252561 91275 253163
rect 86811 252443 91669 252561
rect 91787 252443 91793 252561
rect 86811 252104 86929 252443
rect 90584 252428 90892 252443
rect 86994 252148 87236 252188
rect 86994 252104 87034 252148
rect 86811 251986 87112 252104
rect 85733 251235 85815 251823
rect 86994 251516 87108 251986
rect 87226 251611 87306 252100
rect 87224 251529 87593 251611
rect 87226 251524 87306 251529
rect 86994 251468 87034 251516
rect 86994 251428 87216 251468
rect 86249 251235 86331 251241
rect 87511 251235 87593 251529
rect 85733 251229 87593 251235
rect 85733 251159 86255 251229
rect 86325 251159 87593 251229
rect 85733 251153 87593 251159
rect 86249 251147 86331 251153
rect 86364 250389 86694 251153
rect 86358 250059 86364 250389
rect 86694 250059 86700 250389
rect 87458 241684 87464 242060
rect 87840 241684 87846 242060
rect 87458 241682 87846 241684
rect 81268 238128 85764 239428
rect 79968 238122 81268 238128
rect 79347 235218 83164 235311
rect 83071 232321 83164 235218
rect 84464 235124 85764 238128
rect 84494 232920 85794 233156
rect 87464 232920 87840 241682
rect 111993 239460 112043 270327
rect 118460 269216 118972 269222
rect 118460 268704 118472 269216
rect 118972 268704 118978 269216
rect 118460 268698 118972 268704
rect 123136 243340 123250 330645
rect 204780 307770 219036 307776
rect 124280 299161 131171 299275
rect 131285 299161 131291 299275
rect 124280 243296 124394 299161
rect 202198 298804 204780 307770
rect 202232 295040 204780 298804
rect 170424 293708 204780 295040
rect 170424 293240 199492 293708
rect 199960 293514 204780 293708
rect 219036 302526 219758 307770
rect 219036 293560 219792 302526
rect 199960 293508 219036 293514
rect 199960 293240 206354 293508
rect 125276 267773 131605 267887
rect 131719 267773 131725 267887
rect 125276 243266 125390 267773
rect 170424 264322 171996 293240
rect 199492 293234 199960 293240
rect 215369 291294 215419 291649
rect 209054 291242 209060 291294
rect 209112 291242 209118 291294
rect 215362 291242 215368 291294
rect 215420 291242 215426 291294
rect 209061 290878 209111 291242
rect 209061 290828 209550 290878
rect 211103 290828 211991 290878
rect 211941 290428 211991 290828
rect 211940 290422 211992 290428
rect 211940 290364 211992 290370
rect 224179 290349 225797 362111
rect 582030 300330 582036 300654
rect 582360 300330 582366 300654
rect 582036 299956 582360 300330
rect 581700 299632 582360 299956
rect 581740 296012 581960 299632
rect 579364 295810 579460 295816
rect 578522 295714 579364 295810
rect 579460 295809 579888 295810
rect 579460 295714 579889 295809
rect 581740 295792 582284 296012
rect 578522 294220 578618 295714
rect 579364 295708 579460 295714
rect 581661 295545 581847 295551
rect 581661 295539 581673 295545
rect 579498 295476 579550 295482
rect 579492 295424 579498 295476
rect 579550 295424 579556 295476
rect 579498 295418 579550 295424
rect 581661 295365 581667 295539
rect 581661 295359 581673 295365
rect 581847 295359 581853 295545
rect 581661 295353 581847 295359
rect 579610 295170 579889 295266
rect 581303 295125 581361 295228
rect 581503 295084 581576 295202
rect 582064 295154 582284 295792
rect 581303 295061 581361 295067
rect 581497 295011 581503 295084
rect 581576 295011 581582 295084
rect 581740 294934 582284 295154
rect 579688 294900 579932 294906
rect 581740 294900 581960 294934
rect 579688 294680 579700 294900
rect 579920 294680 581960 294900
rect 579688 294674 579932 294680
rect 579290 294465 580285 294575
rect 579290 294370 579400 294465
rect 578810 294260 579400 294370
rect 580175 294355 580285 294465
rect 579700 294346 579920 294352
rect 578522 294002 578790 294220
rect 578580 290430 578790 294002
rect 578205 290340 578790 290430
rect 578205 290300 578460 290340
rect 578500 290300 578790 290340
rect 578205 290220 578790 290300
rect 579400 294080 579460 294200
rect 580175 294245 580795 294355
rect 579700 294080 579920 294126
rect 580140 294080 580190 294200
rect 579400 290390 580190 294080
rect 579400 290230 579460 290390
rect 580130 290230 580190 290390
rect 580810 294127 581090 294200
rect 580810 294093 581003 294127
rect 581037 294093 581090 294127
rect 580810 294057 581090 294093
rect 581503 294057 581576 294063
rect 580810 293984 581503 294057
rect 580810 293706 581090 293984
rect 581503 293978 581576 293984
rect 580810 293594 583064 293706
rect 583176 293594 583182 293706
rect 580810 290490 581090 293594
rect 581494 290490 581774 290496
rect 577017 289485 577227 289491
rect 578205 289485 578415 290220
rect 580810 290210 581494 290490
rect 581774 290484 582216 290490
rect 581774 290216 581936 290484
rect 582204 290216 582216 290484
rect 581774 290210 582216 290216
rect 581494 290204 581774 290210
rect 578810 290090 579400 290180
rect 580200 290090 580790 290180
rect 579305 289945 579395 290090
rect 580200 289945 580290 290090
rect 579305 289855 583149 289945
rect 579306 289792 583149 289855
rect 579304 289686 583149 289792
rect 580333 289485 580543 289491
rect 577227 289275 580333 289485
rect 580543 289275 581835 289485
rect 577017 289269 577227 289275
rect 580333 289269 580543 289275
rect 199672 282604 200172 282610
rect 214648 282604 215148 288448
rect 217596 287438 225118 288278
rect 573386 287986 573678 287992
rect 573380 287706 573386 287986
rect 573678 287706 573684 287986
rect 573380 287694 573684 287706
rect 164966 263230 171996 264322
rect 164820 263218 171996 263230
rect 164820 262750 165544 263218
rect 166012 262750 171996 263218
rect 174310 282104 199672 282604
rect 200172 282104 215148 282604
rect 164820 262738 165300 262750
rect 163250 262510 163750 262516
rect 174310 262510 174810 282104
rect 199672 282098 200172 282104
rect 217590 279916 217596 287438
rect 225118 279916 225124 287438
rect 163750 262010 174810 262510
rect 581625 275252 581835 289275
rect 581625 275140 581644 275252
rect 581756 275140 581835 275252
rect 163250 262004 163750 262010
rect 165768 257258 166579 257480
rect 166801 257258 168712 257480
rect 168881 256310 168963 256316
rect 168881 256304 168893 256310
rect 168881 256234 168887 256304
rect 168881 256228 168893 256234
rect 168963 256228 168969 256310
rect 168881 256222 168963 256228
rect 168822 256045 168874 256051
rect 168780 255999 168822 256039
rect 168822 255987 168874 255993
rect 165524 255846 165838 255886
rect 165524 249312 165564 255846
rect 167253 255559 167315 255565
rect 167247 255507 167253 255559
rect 167315 255507 167321 255559
rect 167247 255503 167259 255507
rect 167309 255503 167321 255507
rect 167247 255497 167321 255503
rect 168146 254944 168186 255064
rect 168134 254892 168140 254944
rect 168192 254892 168198 254944
rect 195086 253799 195092 254013
rect 195306 253799 195312 254013
rect 166807 253464 166813 253574
rect 166923 253464 166929 253574
rect 167114 252784 167174 253688
rect 167889 253464 167895 253574
rect 168005 253464 168011 253574
rect 167114 252724 170032 252784
rect 165708 250818 166301 251000
rect 166483 250818 168846 251000
rect 169199 249902 169281 249908
rect 169199 249896 169211 249902
rect 169199 249826 169205 249896
rect 169199 249820 169211 249826
rect 169281 249820 169287 249902
rect 169199 249814 169281 249820
rect 169590 249654 169642 249660
rect 168834 249608 169590 249648
rect 169590 249596 169642 249602
rect 161087 249198 165564 249312
rect 126300 244483 126414 244500
rect 126300 244369 131591 244483
rect 131705 244369 131711 244483
rect 126300 243278 126414 244369
rect 161087 241967 161201 249198
rect 165524 249084 165564 249198
rect 165518 249072 165570 249084
rect 165518 249032 165524 249072
rect 165564 249032 165570 249072
rect 165518 249020 165570 249032
rect 167075 248053 167149 248059
rect 167075 248049 167087 248053
rect 167137 248049 167149 248053
rect 167075 247997 167081 248049
rect 167143 247997 167149 248049
rect 167081 247991 167143 247997
rect 169590 247522 169642 247528
rect 166725 247471 166835 247477
rect 169584 247470 169590 247522
rect 169642 247470 169648 247522
rect 169590 247464 169642 247470
rect 166725 247355 166835 247361
rect 167048 246990 167108 247311
rect 167871 247166 167981 247172
rect 167871 247050 167981 247056
rect 169972 246990 170032 252724
rect 162504 246930 170032 246990
rect 161081 241853 161087 241967
rect 161201 241853 161207 241967
rect 119291 239715 119489 239721
rect 119285 239517 119291 239715
rect 119477 239517 119489 239715
rect 119291 239511 119489 239517
rect 111910 239204 112118 239460
rect 111910 238990 112118 238996
rect 123118 237218 123290 237372
rect 124254 237218 124426 237342
rect 125278 237218 125450 237304
rect 126302 237218 126474 237300
rect 123040 236746 126500 237218
rect 121069 235961 121139 235967
rect 121063 235891 121069 235961
rect 121127 235955 121139 235961
rect 121133 235897 121139 235955
rect 121127 235891 121139 235897
rect 121069 235885 121139 235891
rect 89310 235677 89640 235689
rect 89310 235359 89316 235677
rect 89634 235359 89640 235677
rect 89310 235003 89640 235359
rect 89310 232920 89640 234673
rect 124162 234193 124634 236746
rect 161087 234193 161201 241853
rect 124162 234079 161201 234193
rect 84494 232321 91170 232920
rect 83071 232228 91170 232321
rect 84494 231620 91170 232228
rect 92470 231620 92476 232920
rect 84494 231466 85794 231620
rect 124162 230584 124634 234079
rect 162504 232134 162564 246930
rect 163560 246382 164060 246388
rect 163554 245882 163560 246382
rect 164060 245882 164066 246382
rect 166466 246376 166990 246388
rect 163560 245876 164060 245882
rect 166466 245876 166472 246376
rect 166984 245876 166990 246376
rect 166472 245870 166984 245876
rect 173705 245091 173711 245161
rect 173781 245091 173787 245161
rect 173711 245009 173781 245091
rect 181841 244891 181911 244897
rect 181911 244821 183913 244891
rect 181841 244815 181911 244821
rect 163906 243682 164146 243688
rect 163900 243442 163906 243682
rect 164146 243442 164152 243682
rect 163906 243436 164146 243442
rect 128896 232074 129512 232134
rect 129572 232074 162564 232134
rect 124162 230112 159064 230584
rect 84412 228275 85712 229500
rect 124162 228916 124634 230112
rect 124156 228444 124162 228916
rect 124634 228444 124640 228916
rect 84412 228229 85249 228275
rect 85295 228229 85712 228275
rect 84412 227580 85712 228229
rect 84406 226280 84412 227580
rect 85712 226280 85718 227580
rect 158592 206748 159064 230112
rect 168333 223421 168687 223427
rect 168327 223079 168333 223421
rect 168687 223079 168693 223421
rect 168327 223073 168339 223079
rect 168681 223073 168693 223079
rect 168327 223067 168693 223073
rect 159300 220912 159306 221012
rect 159406 220912 174280 221012
rect 174180 220576 174280 220912
rect 175048 220818 175054 220918
rect 175154 220818 175160 220918
rect 177216 220818 177222 220918
rect 177322 220818 177328 220918
rect 175054 220576 175154 220818
rect 174180 220476 175154 220576
rect 177222 220552 177322 220818
rect 195092 220582 195306 253799
rect 581625 237205 581835 275140
rect 582890 269398 583149 289686
rect 582884 269139 582890 269398
rect 583149 269139 583155 269398
rect 581625 236989 581835 236995
rect 197790 221956 208917 222170
rect 209131 221956 209137 222170
rect 197790 220614 198004 221956
rect 177222 220452 185382 220552
rect 173093 220037 173099 220127
rect 173189 220037 175019 220127
rect 183747 219927 185229 220017
rect 183747 216319 183837 219927
rect 183741 216229 183747 216319
rect 183837 216229 183843 216319
rect 194856 213998 198016 214676
rect 194856 213702 198212 213998
rect 175727 209679 175821 212649
rect 185937 210493 186031 212539
rect 185937 210399 192493 210493
rect 192587 210399 192593 210493
rect 175727 209585 192681 209679
rect 192775 209585 192781 209679
rect 197740 206748 198212 213702
rect 158592 206276 198212 206748
<< via1 >>
rect 571508 503354 571560 503366
rect 571508 503320 571514 503354
rect 571514 503320 571554 503354
rect 571554 503320 571560 503354
rect 571508 503314 571560 503320
rect 571482 501586 571630 501588
rect 571482 501440 571626 501586
rect 571626 501440 571630 501586
rect 571482 501438 571630 501440
rect 572150 501414 572342 501606
rect 571516 500775 571568 500784
rect 571516 500741 571525 500775
rect 571525 500741 571559 500775
rect 571559 500741 571568 500775
rect 571516 500732 571568 500741
rect 568903 497307 569053 497457
rect 576654 495826 576898 496070
rect 582222 494146 582282 494206
rect 582142 449278 582845 449981
rect 15182 430948 15762 431528
rect 24690 430264 25750 431324
rect 20362 427598 20822 428058
rect 576272 424294 576372 424394
rect 578922 422439 579097 422614
rect 576630 417764 576742 417876
rect 576580 417651 576703 417657
rect 576580 417540 576586 417651
rect 576586 417540 576697 417651
rect 576697 417540 576703 417651
rect 576580 417534 576703 417540
rect 578953 417729 579479 417735
rect 578953 417215 578959 417729
rect 578959 417215 579473 417729
rect 579473 417215 579479 417729
rect 578953 417209 579479 417215
rect 27813 416171 28663 417021
rect 572822 416070 573022 416270
rect 576324 415982 576376 416034
rect 576324 415122 576376 415174
rect 576324 414880 576376 414932
rect 15937 413887 16591 414541
rect 573594 413340 573646 413392
rect 19894 412852 20016 412974
rect 20302 410761 20512 410971
rect 9304 371169 9546 371411
rect 13980 345166 14040 345172
rect 13980 345118 13986 345166
rect 13986 345118 14034 345166
rect 14034 345118 14040 345166
rect 13980 345112 14040 345118
rect 11826 342944 11878 342950
rect 11826 342904 11832 342944
rect 11832 342904 11872 342944
rect 11872 342904 11878 342944
rect 11826 342898 11878 342904
rect 13485 343601 13567 343607
rect 13485 343537 13491 343601
rect 13491 343537 13561 343601
rect 13561 343537 13567 343601
rect 15499 343589 15617 343595
rect 14087 343567 14139 343573
rect 14087 343517 14133 343567
rect 14133 343517 14139 343567
rect 14087 343511 14139 343517
rect 15499 343483 15505 343589
rect 15505 343483 15611 343589
rect 15611 343483 15617 343589
rect 15499 343477 15617 343483
rect 18117 343471 18235 343601
rect 9262 339834 9494 340066
rect 2248 338350 2636 338356
rect 2248 337980 2254 338350
rect 2254 337980 2630 338350
rect 2630 337980 2636 338350
rect 14314 341306 14366 341358
rect 16397 340623 17247 341473
rect 14740 333562 18584 337406
rect 22866 330765 24484 332383
rect 12111 330581 12233 330691
rect 129751 330645 129865 330759
rect 12244 328276 12512 328544
rect 7492 327840 7544 327892
rect 6128 323962 6588 324422
rect 11773 323988 12623 324838
rect 8336 311186 8440 311290
rect 7492 308794 7544 308846
rect 4892 307618 5482 308208
rect 11708 306280 11908 306480
rect 113634 288820 113734 288920
rect 113448 288280 113548 288380
rect 109990 287510 110042 287562
rect 109126 285798 109626 286298
rect 35044 276629 35182 276767
rect 68793 278362 68894 278463
rect 69939 276404 69993 276458
rect 67455 275949 67561 276055
rect 70495 276404 70549 276458
rect 68547 273645 68657 273755
rect 66047 272603 66849 273405
rect 108900 284224 108952 284276
rect 107588 283874 107640 283926
rect 109470 283814 109522 283866
rect 111114 287498 111166 287550
rect 108226 282104 108278 282156
rect 108470 280018 108522 280070
rect 102999 275869 103129 275999
rect 69825 268339 70439 268603
rect 69825 268250 70087 268339
rect 70087 268250 70176 268339
rect 70176 268250 70439 268339
rect 69825 267989 70439 268250
rect 68261 267361 68591 267691
rect 83334 268345 83948 268603
rect 83334 268244 83591 268345
rect 83591 268244 83692 268345
rect 83692 268244 83948 268345
rect 83334 267989 83948 268244
rect 87108 268500 87244 268636
rect 70836 267156 70968 267288
rect 36697 264895 36790 264988
rect 37439 260287 37532 260380
rect 33483 258839 33553 258909
rect 35564 258712 35616 258764
rect 35778 258712 35830 258764
rect 49864 258744 50020 258900
rect 37508 258434 37592 258518
rect 35448 255144 36082 255778
rect 38630 255178 38734 255282
rect 111330 279020 111382 279072
rect 110595 278415 110765 278421
rect 110595 278245 110759 278415
rect 110759 278245 110765 278415
rect 110595 278239 110765 278245
rect 108979 277437 109153 277489
rect 108979 277399 109075 277437
rect 109075 277399 109113 277437
rect 109113 277399 109153 277437
rect 108979 277315 109153 277399
rect 107811 275869 107941 275999
rect 108534 275778 108586 275830
rect 108534 275046 108586 275098
rect 107562 274328 107614 274380
rect 109466 274268 109518 274320
rect 108080 272933 108132 272985
rect 114920 286880 115400 287348
rect 111620 272574 111720 272580
rect 111620 272486 111626 272574
rect 111626 272486 111714 272574
rect 111714 272486 111720 272574
rect 111620 272480 111720 272486
rect 108424 271070 108476 271122
rect 104884 269296 104988 269400
rect 88653 260629 88983 260959
rect 87447 260504 87505 260510
rect 87447 260446 87499 260504
rect 87499 260446 87505 260504
rect 87447 260440 87505 260446
rect 108424 267274 108924 267280
rect 108424 266786 108430 267274
rect 108430 266786 108918 267274
rect 108918 266786 108924 267274
rect 108424 266780 108924 266786
rect 81153 251203 81159 251307
rect 81159 251203 81269 251307
rect 81269 251203 81275 251307
rect 81153 251197 81275 251203
rect 91365 256693 91417 256699
rect 91365 256643 91371 256693
rect 91371 256643 91417 256693
rect 91365 256637 91417 256643
rect 90584 255694 90892 256002
rect 85345 254623 85519 254797
rect 91669 252443 91787 252561
rect 86364 250059 86694 250389
rect 87464 242052 87840 242060
rect 87464 241688 87470 242052
rect 87470 241688 87834 242052
rect 87834 241688 87840 242052
rect 87464 241684 87840 241688
rect 79968 238128 81268 239428
rect 118472 268704 118972 269216
rect 131171 299161 131285 299275
rect 199492 293240 199960 293708
rect 204780 293514 219036 307770
rect 131605 267773 131719 267887
rect 209060 291242 209112 291294
rect 215368 291242 215420 291294
rect 211940 290370 211992 290422
rect 582036 300330 582360 300654
rect 579364 295714 579460 295810
rect 581673 295539 581847 295545
rect 579498 295470 579550 295476
rect 579498 295430 579504 295470
rect 579504 295430 579544 295470
rect 579544 295430 579550 295470
rect 579498 295424 579550 295430
rect 581673 295365 581841 295539
rect 581841 295365 581847 295539
rect 581673 295359 581847 295365
rect 581303 295067 581361 295125
rect 581503 295011 581576 295084
rect 579700 294680 579920 294900
rect 579700 294126 579920 294346
rect 581503 293984 581576 294057
rect 583064 293594 583176 293706
rect 581494 290210 581774 290490
rect 577017 289275 577227 289485
rect 580333 289275 580543 289485
rect 573386 287706 573678 287986
rect 165544 262750 166012 263218
rect 199672 282104 200172 282604
rect 217596 279916 225118 287438
rect 163250 262010 163750 262510
rect 581644 275140 581756 275252
rect 166579 257258 166801 257480
rect 168893 256304 168963 256310
rect 168893 256234 168957 256304
rect 168957 256234 168963 256304
rect 168893 256228 168963 256234
rect 168822 255993 168874 256045
rect 167253 255553 167315 255559
rect 167253 255507 167259 255553
rect 167259 255507 167309 255553
rect 167309 255507 167315 255553
rect 168140 254892 168192 254944
rect 195092 253799 195306 254013
rect 166813 253568 166923 253574
rect 166813 253470 166819 253568
rect 166819 253470 166917 253568
rect 166917 253470 166923 253568
rect 166813 253464 166923 253470
rect 167895 253464 168005 253574
rect 166301 250818 166483 251000
rect 169211 249896 169281 249902
rect 169211 249826 169275 249896
rect 169275 249826 169281 249896
rect 169211 249820 169281 249826
rect 169590 249602 169642 249654
rect 131591 244369 131705 244483
rect 167081 248003 167087 248049
rect 167087 248003 167137 248049
rect 167137 248003 167143 248049
rect 167081 247997 167143 248003
rect 166725 247361 166835 247471
rect 169590 247516 169642 247522
rect 169590 247476 169596 247516
rect 169596 247476 169636 247516
rect 169636 247476 169642 247516
rect 169590 247470 169642 247476
rect 167871 247056 167981 247166
rect 161087 241853 161201 241967
rect 119291 239517 119477 239715
rect 111910 238996 112118 239204
rect 121069 235955 121127 235961
rect 121069 235897 121075 235955
rect 121075 235897 121127 235955
rect 121069 235891 121127 235897
rect 89310 234673 89640 235003
rect 91170 231620 92470 232920
rect 163560 245882 164060 246382
rect 166472 245876 166984 246376
rect 173711 245091 173781 245161
rect 181841 244821 181911 244891
rect 163906 243442 164146 243682
rect 129512 232074 129572 232134
rect 124162 228444 124634 228916
rect 84412 226280 85712 227580
rect 168333 223415 168687 223421
rect 168333 223079 168339 223415
rect 168339 223079 168681 223415
rect 168681 223079 168687 223415
rect 159306 220912 159406 221012
rect 175054 220818 175154 220918
rect 177222 220818 177322 220918
rect 582890 269139 583149 269398
rect 581625 236995 581835 237205
rect 208917 221956 209131 222170
rect 173099 220037 173189 220127
rect 183747 216229 183837 216319
rect 192493 210399 192587 210493
rect 192681 209585 192775 209679
<< metal2 >>
rect 567957 503522 572531 503765
rect 567957 493513 568200 503522
rect 571508 503366 571560 503372
rect 570955 503323 571508 503357
rect 570955 501035 570989 503323
rect 571508 503308 571560 503314
rect 572288 501606 572531 503522
rect 571462 501588 572150 501606
rect 571462 501438 571482 501588
rect 571630 501438 572150 501588
rect 571462 501414 572150 501438
rect 572342 501414 572976 501606
rect 573168 501414 573177 501606
rect 570955 501001 571559 501035
rect 571525 500784 571559 501001
rect 571510 500732 571516 500784
rect 571568 500732 571574 500784
rect 568903 497457 569053 497463
rect 568894 497307 568903 497457
rect 569053 497307 569062 497457
rect 568903 497301 569053 497307
rect 576654 496070 576898 496076
rect 576645 495826 576654 496070
rect 576898 495826 576907 496070
rect 576654 495820 576898 495826
rect 582213 494146 582222 494206
rect 582282 494146 582291 494206
rect 567957 493270 568672 493513
rect 2340 468340 104146 468452
rect 2340 464869 2452 468340
rect 2336 464767 2345 464869
rect 2447 464767 2456 464869
rect 2340 464762 2452 464767
rect 15182 431528 15762 431534
rect 15173 430948 15182 431528
rect 15762 430948 15771 431528
rect 24690 431324 25750 431330
rect 15182 430942 15762 430948
rect 24681 430264 24690 431324
rect 25750 430264 25759 431324
rect 24690 430258 25750 430264
rect 20362 428058 20822 428064
rect 20353 427598 20362 428058
rect 20822 427598 20831 428058
rect 20362 427592 20822 427598
rect 27818 417021 28658 417025
rect 27807 416171 27813 417021
rect 28663 416171 28669 417021
rect 27818 416167 28658 416171
rect 15931 413887 15937 414541
rect 16591 413887 16597 414541
rect 19894 412974 20016 412983
rect 19888 412852 19894 412974
rect 20016 412852 20022 412974
rect 19894 412843 20016 412852
rect 20302 410971 20512 410977
rect 20293 410761 20302 410971
rect 20512 410761 20521 410971
rect 20302 410755 20512 410761
rect 9304 371411 9546 371417
rect 9295 371169 9304 371411
rect 9546 371169 9555 371411
rect 9304 371163 9546 371169
rect 13434 346865 13704 346874
rect 13434 345476 13704 346595
rect 11813 345336 11822 345396
rect 11882 345336 11891 345396
rect 11832 342950 11872 345336
rect 13491 343607 13561 345476
rect 13982 345396 14038 345403
rect 13980 345394 14040 345396
rect 13980 345338 13982 345394
rect 14038 345338 14040 345394
rect 13980 345172 14040 345338
rect 13974 345112 13980 345172
rect 14040 345112 14046 345172
rect 13479 343537 13485 343607
rect 13567 343537 13573 343607
rect 18117 343601 18235 343607
rect 14087 343573 14139 343579
rect 14074 343511 14083 343573
rect 14143 343511 14152 343573
rect 14087 343505 14139 343511
rect 15493 343477 15499 343595
rect 15617 343477 18117 343595
rect 18235 343471 18237 343595
rect 18117 343465 18237 343471
rect 11820 342898 11826 342950
rect 11878 342898 11884 342950
rect 11832 341048 11872 342898
rect 16397 341473 17247 341479
rect 14310 341362 14370 341371
rect 14308 341306 14310 341358
rect 14370 341306 14372 341358
rect 14310 341293 14370 341302
rect 2850 340588 11872 341048
rect 16393 340628 16397 341468
rect 17247 340628 17251 341468
rect 16397 340617 17247 340623
rect 2248 338356 2636 338365
rect 2242 337980 2248 338356
rect 2636 337980 2642 338356
rect 2248 337971 2636 337980
rect 2850 324422 3310 340588
rect 9262 340066 9494 340075
rect 9256 339834 9262 340066
rect 9494 339834 9500 340066
rect 9262 339825 9494 339834
rect 18119 338566 18237 343465
rect 18024 338258 90892 338566
rect 14740 337406 18584 337412
rect 14731 333562 14740 337406
rect 18584 333562 18593 337406
rect 14740 333556 18584 333562
rect 22866 332383 24484 332389
rect 22862 330770 22866 332378
rect 24484 330770 24488 332378
rect 22866 330759 24484 330765
rect 12111 330691 12233 330700
rect 12105 330581 12111 330691
rect 12233 330581 12239 330691
rect 12111 330572 12233 330581
rect 12244 328544 12512 328550
rect 12235 328276 12244 328544
rect 12512 328276 12521 328544
rect 12244 328270 12512 328276
rect 7486 327840 7492 327892
rect 7544 327840 7550 327892
rect 6128 324422 6588 324428
rect 2850 323962 6128 324422
rect 6128 323956 6588 323962
rect 7493 308846 7543 327840
rect 11773 324838 12623 324847
rect 11767 323988 11773 324838
rect 12623 323988 12629 324838
rect 11773 323979 12623 323988
rect 8336 311290 8440 311296
rect 8332 311191 8336 311285
rect 8440 311191 8444 311285
rect 8336 311180 8440 311186
rect 7486 308794 7492 308846
rect 7544 308794 7550 308846
rect 4892 308208 5482 308217
rect 4886 307618 4892 308208
rect 5482 307618 5488 308208
rect 4892 307609 5482 307618
rect 11708 306480 11908 306486
rect 11699 306280 11708 306480
rect 11908 306280 11917 306480
rect 11708 306274 11908 306280
rect 2717 300636 2726 301936
rect 4026 300636 4035 301936
rect 2726 236469 4026 300636
rect 9200 292860 10500 292869
rect 5348 291560 9200 292860
rect 2722 235179 2731 236469
rect 4021 235179 4030 236469
rect 2726 235174 4026 235179
rect 5348 227575 6648 291560
rect 9200 291551 10500 291560
rect 68793 278463 68894 278472
rect 68787 278362 68793 278463
rect 68894 278362 68900 278463
rect 68793 278353 68894 278362
rect 35044 276767 35182 276773
rect 35035 276629 35044 276767
rect 35182 276629 35191 276767
rect 35044 276623 35182 276629
rect 69933 276404 69939 276458
rect 69993 276404 70495 276458
rect 70549 276404 70555 276458
rect 67455 276055 67561 276061
rect 67446 275949 67455 276055
rect 67561 275949 67570 276055
rect 67455 275943 67561 275949
rect 68547 273755 68657 273764
rect 68541 273645 68547 273755
rect 68657 273645 68663 273755
rect 68547 273636 68657 273645
rect 66052 273405 66844 273409
rect 66041 272603 66047 273405
rect 66849 272603 66855 273405
rect 66052 272599 66844 272603
rect 37670 268584 40976 268668
rect 41060 268584 41069 268668
rect 87108 268636 87244 268645
rect 69825 268603 70439 268609
rect 83334 268603 83948 268609
rect 36697 264988 36790 264994
rect 36688 264895 36697 264988
rect 36790 264895 36799 264988
rect 36697 264889 36790 264895
rect 37439 260380 37532 260386
rect 37430 260287 37439 260380
rect 37532 260287 37541 260380
rect 37439 260281 37532 260287
rect 37670 259892 37754 268584
rect 69821 267994 69825 268598
rect 70439 267994 70443 268598
rect 83325 267989 83334 268603
rect 83948 267989 83957 268603
rect 87102 268500 87108 268636
rect 87244 268500 87250 268636
rect 87108 268491 87244 268500
rect 69825 267983 70439 267989
rect 83334 267983 83948 267989
rect 68261 267691 68591 267697
rect 68257 267366 68261 267686
rect 68591 267366 68595 267686
rect 68261 267355 68591 267361
rect 70836 267288 70968 267297
rect 70830 267156 70836 267288
rect 70968 267156 70974 267288
rect 70836 267147 70968 267156
rect 88658 260959 88978 260963
rect 88647 260629 88653 260959
rect 88983 260629 88989 260959
rect 88658 260625 88978 260629
rect 87447 260510 87505 260516
rect 87437 260440 87446 260510
rect 87506 260440 87515 260510
rect 87447 260434 87505 260440
rect 37508 259808 37754 259892
rect 33483 258909 33553 258918
rect 33483 258830 33553 258839
rect 35564 258764 35616 258770
rect 35772 258758 35778 258764
rect 35616 258718 35778 258758
rect 35772 258712 35778 258718
rect 35830 258712 35836 258764
rect 35564 258706 35616 258712
rect 37508 258518 37592 259808
rect 49864 258900 50020 258906
rect 49855 258744 49864 258900
rect 50020 258744 50029 258900
rect 49864 258738 50020 258744
rect 37502 258434 37508 258518
rect 37592 258434 37598 258518
rect 90584 257328 90892 338258
rect 104034 289130 104146 468340
rect 568429 412864 568672 493270
rect 582142 449981 582845 449987
rect 582133 449278 582142 449981
rect 582845 449278 582854 449981
rect 582142 449272 582845 449278
rect 576272 424394 576372 424400
rect 576263 424294 576272 424394
rect 576372 424294 576381 424394
rect 576272 424288 576372 424294
rect 578922 422614 579097 422620
rect 578913 422439 578922 422614
rect 579097 422439 579106 422614
rect 578922 422433 579097 422439
rect 576635 417876 576737 417880
rect 576624 417764 576630 417876
rect 576742 417764 576748 417876
rect 576635 417760 576737 417764
rect 578953 417735 579479 417741
rect 576289 417534 576580 417657
rect 576703 417534 576709 417657
rect 576289 416467 576412 417534
rect 578949 417214 578953 417730
rect 579479 417214 579483 417730
rect 578953 417203 579479 417209
rect 572822 416270 573022 416279
rect 572816 416070 572822 416270
rect 573022 416070 573028 416270
rect 572822 416061 573022 416070
rect 576326 416034 576374 416467
rect 576318 415982 576324 416034
rect 576376 415982 576382 416034
rect 575985 415780 577187 415930
rect 576324 415174 576376 415180
rect 576324 415116 576376 415122
rect 576326 414932 576374 415116
rect 576318 414880 576324 414932
rect 576376 414880 576382 414932
rect 577037 414665 577187 415780
rect 577037 414515 578359 414665
rect 578509 414515 578518 414665
rect 573588 413340 573594 413392
rect 573646 413340 573652 413392
rect 573597 412864 573643 413340
rect 568429 412621 573742 412864
rect 129751 330759 129865 330765
rect 129742 330645 129751 330759
rect 129865 330645 129874 330759
rect 129751 330639 129865 330645
rect 155850 323300 156002 323309
rect 156002 323249 156372 323300
rect 156002 323199 167309 323249
rect 156002 323148 156372 323199
rect 155850 323139 156002 323148
rect 128168 305774 128224 305781
rect 128166 305772 128226 305774
rect 128166 305716 128168 305772
rect 128224 305716 128226 305772
rect 128166 300898 128226 305716
rect 104032 289018 104146 289130
rect 104034 288632 104146 289018
rect 123612 300838 128226 300898
rect 113634 288920 113734 288926
rect 113625 288820 113634 288920
rect 113734 288820 113743 288920
rect 113634 288814 113734 288820
rect 104032 288520 104434 288632
rect 113448 288380 113548 288386
rect 113439 288280 113448 288380
rect 113548 288280 113557 288380
rect 113448 288274 113548 288280
rect 109991 287568 110041 288235
rect 110525 287683 110575 288213
rect 110525 287633 110951 287683
rect 109990 287562 110042 287568
rect 109990 287504 110042 287510
rect 109126 286298 109626 286304
rect 109122 285803 109126 286293
rect 109626 285803 109630 286293
rect 109126 285792 109626 285798
rect 108901 285346 108951 285390
rect 110148 285346 110204 285353
rect 108901 285344 110206 285346
rect 108901 285288 110148 285344
rect 110204 285288 110206 285344
rect 108901 285286 110206 285288
rect 108901 284282 108951 285286
rect 110148 285279 110204 285286
rect 108900 284276 108952 284282
rect 108900 284218 108952 284224
rect 107584 283930 107644 283939
rect 107582 283874 107584 283926
rect 107644 283874 107646 283926
rect 109470 283870 109522 283872
rect 107584 283861 107644 283870
rect 109457 283810 109466 283870
rect 109526 283810 109535 283870
rect 109470 283808 109522 283810
rect 108226 282156 108278 282162
rect 110901 282155 110951 287633
rect 111115 287550 111165 288201
rect 111703 287715 111753 288245
rect 111703 287665 112795 287715
rect 111108 287498 111114 287550
rect 111166 287498 111172 287550
rect 111292 285006 111352 285008
rect 111285 284950 111294 285006
rect 111350 284950 111359 285006
rect 111292 283586 111352 284950
rect 111292 283520 111381 283586
rect 108278 282105 110951 282155
rect 108226 282098 108278 282104
rect 108464 280018 108470 280070
rect 108522 280018 108528 280070
rect 108471 277967 108521 280018
rect 111331 279072 111381 283520
rect 111324 279020 111330 279072
rect 111382 279020 111388 279072
rect 110595 278421 110765 278427
rect 110586 278239 110595 278421
rect 110765 278239 110774 278421
rect 110595 278233 110765 278239
rect 110396 277967 110496 277992
rect 108471 277917 110496 277967
rect 110396 277726 110496 277917
rect 110387 277626 110396 277726
rect 110496 277626 110505 277726
rect 108979 277489 109153 277495
rect 102427 277315 108979 277489
rect 102427 266679 102601 277315
rect 108979 277309 109153 277315
rect 102999 275999 103129 276005
rect 107811 275999 107941 276005
rect 103129 275869 107811 275999
rect 102999 275863 103129 275869
rect 107811 275863 107941 275869
rect 108528 275778 108534 275830
rect 108586 275778 108592 275830
rect 108535 275098 108585 275778
rect 108528 275046 108534 275098
rect 108586 275046 108592 275098
rect 107562 274384 107614 274386
rect 107549 274324 107558 274384
rect 107618 274324 107627 274384
rect 109466 274324 109518 274326
rect 107562 274322 107614 274324
rect 109453 274264 109462 274324
rect 109522 274264 109531 274324
rect 109466 274262 109518 274264
rect 108074 272933 108080 272985
rect 108132 272933 108138 272985
rect 108081 272880 108131 272933
rect 108081 272869 108137 272880
rect 112745 272869 112795 287665
rect 114920 287348 115400 287357
rect 114914 286880 114920 287348
rect 115400 286880 115406 287348
rect 114920 286871 115400 286880
rect 113783 283974 113792 284034
rect 113852 283974 113861 284034
rect 113792 282692 113852 283974
rect 123612 282692 123672 300838
rect 131171 299275 131285 299281
rect 131162 299161 131171 299275
rect 131285 299161 131294 299275
rect 131171 299155 131285 299161
rect 113792 282632 123672 282692
rect 108081 272841 112795 272869
rect 108087 272819 112795 272841
rect 111620 272580 111720 272586
rect 111620 272034 111720 272480
rect 109756 271934 111720 272034
rect 108424 271122 108476 271128
rect 108476 271071 108681 271121
rect 108424 271064 108476 271070
rect 104884 269400 104988 269406
rect 104880 269301 104884 269395
rect 104988 269301 104992 269395
rect 104884 269290 104988 269296
rect 108631 267286 108681 271071
rect 108424 267280 108924 267286
rect 108420 266785 108424 267275
rect 108924 266785 108928 267275
rect 109756 267252 109856 271934
rect 118472 269216 118972 269222
rect 119831 269210 120321 269212
rect 118972 269203 125164 269210
rect 118972 268713 119831 269203
rect 120321 268713 125164 269203
rect 118972 268710 125164 268713
rect 119826 268708 122388 268710
rect 119831 268704 120321 268708
rect 118472 268698 118972 268704
rect 109756 267152 120556 267252
rect 108424 266774 108924 266780
rect 90584 257011 90892 257020
rect 91327 266505 102601 266679
rect 91327 256735 91501 266505
rect 120456 258908 120556 267152
rect 124664 262510 125164 268710
rect 131605 267887 131719 267893
rect 131596 267773 131605 267887
rect 131719 267773 131728 267887
rect 131605 267767 131719 267773
rect 157327 264306 157525 264315
rect 157525 264215 158346 264306
rect 157525 264165 164553 264215
rect 157525 264108 158346 264165
rect 157327 264099 157525 264108
rect 124664 262010 163250 262510
rect 163750 262010 164060 262510
rect 120456 258808 129026 258908
rect 84749 256699 91501 256735
rect 84749 256637 91365 256699
rect 91417 256637 91501 256699
rect 84749 256561 91501 256637
rect 84749 256524 84923 256561
rect 84745 256360 84754 256524
rect 84918 256360 84927 256524
rect 84749 256355 84923 256360
rect 90584 256002 90892 256008
rect 35448 255778 36082 255787
rect 35442 255144 35448 255778
rect 36082 255144 36088 255778
rect 90580 255699 90584 255997
rect 90892 255699 90896 255997
rect 90584 255688 90892 255694
rect 38635 255282 38729 255286
rect 38624 255178 38630 255282
rect 38734 255178 38740 255282
rect 38635 255174 38729 255178
rect 35448 255135 36082 255144
rect 85345 254797 85519 254803
rect 85336 254623 85345 254797
rect 85519 254623 85528 254797
rect 85345 254617 85519 254623
rect 91669 252561 91787 252567
rect 91660 252443 91669 252561
rect 91787 252443 91796 252561
rect 91669 252437 91787 252443
rect 81153 251307 81275 251316
rect 81147 251197 81153 251307
rect 81275 251197 81281 251307
rect 81153 251188 81275 251197
rect 86364 250389 86694 250395
rect 86355 250059 86364 250389
rect 86694 250059 86703 250389
rect 86364 250053 86694 250059
rect 87464 242060 87840 242066
rect 87455 241684 87464 242060
rect 87840 241684 87849 242060
rect 87464 241678 87840 241684
rect 119291 239715 119477 239721
rect 119282 239517 119291 239715
rect 119477 239602 119486 239715
rect 119477 239542 119954 239602
rect 119477 239517 119486 239542
rect 119291 239511 119477 239517
rect 79968 239428 81268 239437
rect 79962 238128 79968 239428
rect 81268 238128 81274 239428
rect 111910 239204 112118 239213
rect 111904 238996 111910 239204
rect 112118 238996 112124 239204
rect 111910 238987 112118 238996
rect 79968 238119 81268 238128
rect 89310 235003 89640 235012
rect 89304 234673 89310 235003
rect 89640 234673 89646 235003
rect 89310 234664 89640 234673
rect 91170 232920 92470 232926
rect 91161 231620 91170 232920
rect 92470 231620 92479 232920
rect 119894 232134 119954 239542
rect 121069 235961 121127 235967
rect 121059 235891 121068 235961
rect 121128 235891 121137 235961
rect 121069 235885 121127 235891
rect 128926 234962 129026 258808
rect 163560 246452 164060 262010
rect 164503 248387 164553 264165
rect 165544 263218 166012 263224
rect 165535 262750 165544 263218
rect 166012 262750 166021 263218
rect 165544 262744 166012 262750
rect 166579 257480 166801 257486
rect 166570 257258 166579 257480
rect 166801 257258 166810 257480
rect 166579 257252 166801 257258
rect 167259 255559 167309 323199
rect 204780 307770 219036 307779
rect 199492 293708 199960 293717
rect 199486 293240 199492 293708
rect 199960 293240 199966 293708
rect 204774 293514 204780 307770
rect 219036 293514 219042 307770
rect 582036 300654 582360 300660
rect 582032 300335 582036 300649
rect 582360 300335 582364 300649
rect 582036 300324 582360 300330
rect 579364 295810 579460 295819
rect 579358 295714 579364 295810
rect 579460 295714 579466 295810
rect 579364 295705 579460 295714
rect 581673 295545 581847 295551
rect 579492 295424 579498 295476
rect 579550 295424 579556 295476
rect 579504 294768 579544 295424
rect 581664 295359 581673 295545
rect 581847 295359 581856 295545
rect 581673 295353 581847 295359
rect 581293 295066 581302 295126
rect 581362 295066 581371 295126
rect 581503 295084 581576 295090
rect 579700 294900 579920 294906
rect 579504 294728 579700 294768
rect 579700 294346 579920 294680
rect 579694 294126 579700 294346
rect 579920 294126 579926 294346
rect 581503 294057 581576 295011
rect 581497 293984 581503 294057
rect 581576 293984 581582 294057
rect 583064 293706 583176 293712
rect 583060 293599 583064 293701
rect 583176 293599 583180 293701
rect 583064 293588 583176 293594
rect 204780 293505 219036 293514
rect 199492 293231 199960 293240
rect 209060 291294 209112 291300
rect 215368 291294 215420 291300
rect 209112 291243 215368 291293
rect 209060 291236 209112 291242
rect 215368 291236 215420 291242
rect 581494 290490 581774 290499
rect 211934 290370 211940 290422
rect 211992 290370 211998 290422
rect 199672 282604 200172 282613
rect 199666 282104 199672 282604
rect 200172 282104 200178 282604
rect 199672 282095 200172 282104
rect 211941 274928 211991 290370
rect 581488 290210 581494 290490
rect 581774 290210 581780 290490
rect 581494 290201 581774 290210
rect 577017 289485 577227 289494
rect 580333 289485 580543 289494
rect 577011 289275 577017 289485
rect 577227 289275 577233 289485
rect 580327 289275 580333 289485
rect 580543 289275 580549 289485
rect 577017 289266 577227 289275
rect 580333 289266 580543 289275
rect 573386 287986 573678 287995
rect 573380 287706 573386 287986
rect 573678 287706 573684 287986
rect 573386 287697 573678 287706
rect 217596 287438 225118 287444
rect 217587 279916 217596 287438
rect 225118 279916 225127 287438
rect 217596 279910 225118 279916
rect 581644 275252 581756 275258
rect 581640 275145 581644 275247
rect 581756 275145 581760 275247
rect 581644 275134 581756 275140
rect 211911 274817 213030 274928
rect 213141 274817 213150 274928
rect 582890 269398 583149 269404
rect 582881 269139 582890 269398
rect 583149 269139 583158 269398
rect 582890 269133 583149 269139
rect 168893 256310 168963 256316
rect 168963 256234 169943 256304
rect 168893 256222 168963 256228
rect 168816 255993 168822 256045
rect 168874 255993 168880 256045
rect 167247 255507 167253 255559
rect 167315 255507 167321 255559
rect 168828 255326 168868 255993
rect 169095 255326 169236 255330
rect 168828 255321 169241 255326
rect 168828 255180 169095 255321
rect 169236 255180 169241 255321
rect 168828 255175 169241 255180
rect 168140 254944 168192 254950
rect 168828 254938 168868 255175
rect 169095 255171 169236 255175
rect 168192 254898 168868 254938
rect 168140 254886 168192 254892
rect 166813 253574 166923 253580
rect 167895 253574 168005 253580
rect 166923 253464 167895 253574
rect 166813 253458 166923 253464
rect 167337 253169 167447 253464
rect 167895 253458 168005 253464
rect 167328 253059 167337 253169
rect 167447 253059 167456 253169
rect 166301 251000 166483 251006
rect 166292 250818 166301 251000
rect 166483 250818 166492 251000
rect 166301 250812 166483 250818
rect 169873 250311 169943 256234
rect 195092 254013 195306 254019
rect 195083 253799 195092 254013
rect 195306 253799 195315 254013
rect 195092 253793 195306 253799
rect 169873 250241 172941 250311
rect 169211 249902 169281 249908
rect 169281 249826 170971 249896
rect 169211 249814 169281 249820
rect 169584 249602 169590 249654
rect 169642 249602 169648 249654
rect 164503 248337 167137 248387
rect 167087 248049 167137 248337
rect 167075 247997 167081 248049
rect 167143 247997 167149 248049
rect 169596 247522 169636 249602
rect 166719 247361 166725 247471
rect 166835 247361 166841 247471
rect 169584 247470 169590 247522
rect 169642 247470 169648 247522
rect 166725 246452 166835 247361
rect 167865 247056 167871 247166
rect 167981 247056 167987 247166
rect 163560 246385 166976 246452
rect 163560 246382 166984 246385
rect 163554 245882 163560 246382
rect 164060 246376 166984 246382
rect 164060 245952 166472 246376
rect 164060 245882 164066 245952
rect 166466 245876 166472 245952
rect 166984 246251 166990 246376
rect 167871 246251 167981 247056
rect 166984 246141 167981 246251
rect 166984 245876 166990 246141
rect 166472 245867 166984 245876
rect 159711 245292 159720 245428
rect 159856 245390 160634 245428
rect 169596 245390 169636 247470
rect 159856 245350 169636 245390
rect 159856 245292 160634 245350
rect 170901 245161 170971 249826
rect 172871 246537 172941 250241
rect 172871 246467 181911 246537
rect 173711 245161 173781 245167
rect 170901 245091 173711 245161
rect 173711 245085 173781 245091
rect 181841 244891 181911 246467
rect 181835 244821 181841 244891
rect 181911 244821 181917 244891
rect 131591 244483 131705 244489
rect 131582 244369 131591 244483
rect 131705 244369 131714 244483
rect 131591 244363 131705 244369
rect 163906 243682 164146 243688
rect 163902 243447 163906 243677
rect 164146 243447 164150 243677
rect 163906 243436 164146 243442
rect 161087 241967 161201 241973
rect 161078 241853 161087 241967
rect 161201 241853 161210 241967
rect 161087 241847 161201 241853
rect 161573 237279 161855 237288
rect 161855 236997 165169 237279
rect 161573 236988 161855 236997
rect 128926 234862 145650 234962
rect 129512 232134 129572 232140
rect 119894 232074 129512 232134
rect 129512 232068 129572 232074
rect 91170 231614 92470 231620
rect 124162 228916 124634 228922
rect 124153 228444 124162 228916
rect 124634 228444 124643 228916
rect 124162 228438 124634 228444
rect 84412 227580 85712 227586
rect 5348 226285 5353 227575
rect 6643 226285 6648 227575
rect 5348 226280 6648 226285
rect 84403 226280 84412 227580
rect 85712 226280 85721 227580
rect 5353 226276 6643 226280
rect 84412 226274 85712 226280
rect 145550 221012 145650 234862
rect 159306 221012 159406 221018
rect 145550 220912 159306 221012
rect 159306 220906 159406 220912
rect 164887 220405 165169 236997
rect 581616 236995 581625 237205
rect 581835 236995 581844 237205
rect 168333 223421 168687 223430
rect 168327 223079 168333 223421
rect 168687 223079 168693 223421
rect 168333 223070 168687 223079
rect 208917 222170 209131 222176
rect 208908 221956 208917 222170
rect 209131 221956 209140 222170
rect 208917 221950 209131 221956
rect 175054 220918 175154 220924
rect 177222 220918 177322 220924
rect 175154 220818 177222 220918
rect 175054 220812 175154 220818
rect 177222 220812 177322 220818
rect 172036 220405 172318 220410
rect 164887 220127 172318 220405
rect 173099 220127 173189 220133
rect 164887 220123 173099 220127
rect 164887 198319 165169 220123
rect 172036 220037 173099 220123
rect 172036 219872 172318 220037
rect 173099 220031 173189 220037
rect 172223 216319 172313 219872
rect 183747 216319 183837 216325
rect 172223 216229 183747 216319
rect 183747 216223 183837 216229
rect 192493 210493 192587 210499
rect 192484 210399 192493 210493
rect 192587 210399 192596 210493
rect 192493 210393 192587 210399
rect 192681 209679 192775 209685
rect 192672 209585 192681 209679
rect 192775 209585 192784 209679
rect 192681 209579 192775 209585
rect 164878 198037 164887 198319
rect 165169 198037 165178 198319
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 572976 501414 573168 501606
rect 568903 497307 569053 497457
rect 576654 495826 576898 496070
rect 582222 494146 582282 494206
rect 2345 464767 2447 464869
rect 15182 430948 15762 431528
rect 24690 430264 25750 431324
rect 20362 427598 20822 428058
rect 27818 416176 28658 417016
rect 15942 413892 16586 414536
rect 19894 412852 20016 412974
rect 20302 410761 20512 410971
rect 9304 371169 9546 371411
rect 13434 346595 13704 346865
rect 11822 345336 11882 345396
rect 13982 345338 14038 345394
rect 14083 343511 14087 343573
rect 14087 343511 14139 343573
rect 14139 343511 14143 343573
rect 14310 341358 14370 341362
rect 14310 341306 14314 341358
rect 14314 341306 14366 341358
rect 14366 341306 14370 341358
rect 14310 341302 14370 341306
rect 16402 340628 17242 341468
rect 2248 337980 2636 338356
rect 9262 339834 9494 340066
rect 14740 333562 18584 337406
rect 22871 330770 24479 332378
rect 12111 330581 12233 330691
rect 12244 328276 12512 328544
rect 11773 323988 12623 324838
rect 8341 311191 8435 311285
rect 4892 307618 5482 308208
rect 11708 306280 11908 306480
rect 2726 300636 4026 301936
rect 9200 291560 10500 292860
rect 2731 235179 4021 236469
rect 68793 278362 68894 278463
rect 35044 276629 35182 276767
rect 67455 275949 67561 276055
rect 68547 273645 68657 273755
rect 66052 272608 66844 273400
rect 40976 268584 41060 268668
rect 36697 264895 36790 264988
rect 37439 260287 37532 260380
rect 69830 267994 70434 268598
rect 83334 267989 83948 268603
rect 87108 268500 87244 268636
rect 68266 267366 68586 267686
rect 70836 267156 70968 267288
rect 88658 260634 88978 260954
rect 87446 260440 87447 260510
rect 87447 260440 87505 260510
rect 87505 260440 87506 260510
rect 33483 258839 33553 258909
rect 49864 258744 50020 258900
rect 582142 449278 582845 449981
rect 576272 424294 576372 424394
rect 578922 422439 579097 422614
rect 576635 417769 576737 417871
rect 578958 417214 579474 417730
rect 572822 416070 573022 416270
rect 578359 414515 578509 414665
rect 129751 330645 129865 330759
rect 155850 323148 156002 323300
rect 128168 305716 128224 305772
rect 113634 288820 113734 288920
rect 113448 288280 113548 288380
rect 109131 285803 109621 286293
rect 110148 285288 110204 285344
rect 107584 283926 107644 283930
rect 107584 283874 107588 283926
rect 107588 283874 107640 283926
rect 107640 283874 107644 283926
rect 107584 283870 107644 283874
rect 109466 283866 109526 283870
rect 109466 283814 109470 283866
rect 109470 283814 109522 283866
rect 109522 283814 109526 283866
rect 109466 283810 109526 283814
rect 111294 284950 111350 285006
rect 110595 278239 110765 278421
rect 110396 277626 110496 277726
rect 107558 274380 107618 274384
rect 107558 274328 107562 274380
rect 107562 274328 107614 274380
rect 107614 274328 107618 274380
rect 107558 274324 107618 274328
rect 109462 274320 109522 274324
rect 109462 274268 109466 274320
rect 109466 274268 109518 274320
rect 109518 274268 109522 274320
rect 109462 274264 109522 274268
rect 114920 286880 115400 287348
rect 113792 283974 113852 284034
rect 131171 299161 131285 299275
rect 104889 269301 104983 269395
rect 108429 266785 108919 267275
rect 119831 268713 120321 269203
rect 90584 257020 90892 257328
rect 131605 267773 131719 267887
rect 157327 264108 157525 264306
rect 84754 256360 84918 256524
rect 35448 255144 36082 255778
rect 90589 255699 90887 255997
rect 38635 255183 38729 255277
rect 85345 254623 85519 254797
rect 91669 252443 91787 252561
rect 81153 251197 81275 251307
rect 86364 250059 86694 250389
rect 87464 241684 87840 242060
rect 119291 239517 119477 239715
rect 79968 238128 81268 239428
rect 111910 238996 112118 239204
rect 89310 234673 89640 235003
rect 91170 231620 92470 232920
rect 121068 235891 121069 235961
rect 121069 235891 121127 235961
rect 121127 235891 121128 235961
rect 165544 262750 166012 263218
rect 166579 257258 166801 257480
rect 199492 293240 199960 293708
rect 204780 293514 219036 307770
rect 582041 300335 582355 300649
rect 579364 295714 579460 295810
rect 581673 295359 581847 295545
rect 581302 295125 581362 295126
rect 581302 295067 581303 295125
rect 581303 295067 581361 295125
rect 581361 295067 581362 295125
rect 581302 295066 581362 295067
rect 583069 293599 583171 293701
rect 199672 282104 200172 282604
rect 581494 290210 581774 290490
rect 577017 289275 577227 289485
rect 580333 289275 580543 289485
rect 573386 287706 573678 287986
rect 217596 279916 225118 287438
rect 581649 275145 581751 275247
rect 213030 274817 213141 274928
rect 582890 269139 583149 269398
rect 169095 255180 169236 255321
rect 167337 253059 167447 253169
rect 166301 250818 166483 251000
rect 195092 253799 195306 254013
rect 166472 245876 166984 246376
rect 159720 245292 159856 245428
rect 131591 244369 131705 244483
rect 163911 243447 164141 243677
rect 161087 241853 161201 241967
rect 161573 236997 161855 237279
rect 124162 228444 124634 228916
rect 5353 226285 6643 227575
rect 84412 226280 85712 227580
rect 581625 236995 581835 237205
rect 168333 223079 168687 223421
rect 208917 221956 209131 222170
rect 192493 210399 192587 210493
rect 192681 209585 192775 209679
rect 164887 198037 165169 198319
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702300 73194 704800
rect 120194 702300 125194 704800
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 702300 418394 704800
rect 465394 702300 470394 704800
rect 510594 702340 515394 704800
rect 520594 702340 525394 704800
rect 566594 702300 571594 704800
rect -800 680242 1700 685242
rect 582300 677984 584800 682984
rect -800 643842 1660 648642
rect 582340 639784 584800 644584
rect -800 633842 1660 638642
rect 582340 629784 584800 634584
rect 583004 589584 583116 589590
rect 583116 589472 583234 589584
rect 583004 589466 583116 589472
rect 583356 589472 584800 589584
rect 581842 588520 582251 588529
rect 573686 588420 582251 588520
rect 573686 588402 582412 588420
rect 573686 588290 584800 588402
rect 573686 588228 582412 588290
rect 573686 587146 582251 588228
rect 573686 587060 581988 587146
rect 583520 587108 584800 587220
rect -800 559442 1660 564242
rect -800 549442 1660 554242
rect -800 511530 480 511642
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect 572971 501606 573173 501611
rect 573686 501606 575146 587060
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 583520 583562 584800 583674
rect 582340 550562 584800 555362
rect 582340 540562 584800 545362
rect 572971 501414 572976 501606
rect 573168 501452 575146 501606
rect 573168 501414 573876 501452
rect 572971 501409 573173 501414
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 568892 497302 568898 497462
rect 569048 497457 569058 497462
rect 569053 497307 569058 497457
rect 569048 497302 569058 497307
rect 583520 496504 584800 496616
rect 576649 496070 576659 496075
rect 576649 495826 576654 496070
rect 576649 495821 576659 495826
rect 576903 495821 576909 496075
rect 583520 495322 584800 495434
rect 582217 494206 582287 494211
rect 583520 494206 584800 494252
rect 582217 494146 582222 494206
rect 582282 494146 584800 494206
rect 582217 494141 582287 494146
rect 583520 494140 584800 494146
rect 576194 485746 578654 488408
rect 579365 485746 581823 485751
rect 576194 485745 581824 485746
rect 576194 483287 579365 485745
rect 581823 483287 581824 485745
rect 576194 483286 581824 483287
rect 579365 483281 581823 483286
rect -800 468308 480 468420
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464869 2452 464874
rect -800 464767 2345 464869
rect 2447 464767 2452 464869
rect -800 464762 2452 464767
rect -800 463580 480 463692
rect 18616 462510 18728 462516
rect -800 462398 12902 462510
rect 13008 462398 18616 462510
rect 18616 462392 18728 462398
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 578044 448099 580504 452832
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 582137 449981 582850 449986
rect 582137 449278 582142 449981
rect 582845 449808 583257 449981
rect 583520 449808 584800 449830
rect 582845 449720 584800 449808
rect 582845 449278 583257 449720
rect 583520 449718 584800 449720
rect 582137 449273 582850 449278
rect 578044 448094 581823 448099
rect 578044 448093 581824 448094
rect 578044 445635 579365 448093
rect 581823 445635 581824 448093
rect 578044 445634 581824 445635
rect 579365 445629 581823 445634
rect 15177 431528 15187 431533
rect 15177 430948 15182 431528
rect 15177 430943 15187 430948
rect 15767 430943 15773 431533
rect 24685 431324 25755 431329
rect 21372 430264 24690 431324
rect 25750 430264 25755 431324
rect 24685 430259 25755 430264
rect 20357 428058 20827 428063
rect 1788 427598 20362 428058
rect 20822 427598 20827 428058
rect 1788 425376 2248 427598
rect 20357 427593 20827 427598
rect 992 425198 2248 425376
rect -800 425086 2248 425198
rect 992 424916 2248 425086
rect 576261 424289 576267 424399
rect 576367 424394 576377 424399
rect 576372 424294 576377 424394
rect 576367 424289 576377 424294
rect -800 423904 480 424016
rect -800 422722 480 422834
rect 578917 422614 578927 422619
rect 578917 422439 578922 422614
rect 578917 422434 578927 422439
rect 579102 422434 579108 422619
rect -800 421540 480 421652
rect -800 420358 480 420470
rect -800 419176 480 419288
rect 576630 417871 576940 417876
rect 576630 417769 576635 417871
rect 576737 417769 576940 417871
rect 576630 417764 576940 417769
rect 27814 417021 28662 417026
rect 27813 417020 28663 417021
rect 27813 416172 27814 417020
rect 28662 416172 28663 417020
rect 27813 416171 28663 416172
rect 572817 416275 573027 416281
rect 27814 416166 28662 416171
rect 572817 416070 572822 416075
rect 573022 416070 573027 416075
rect 572817 416065 573027 416070
rect 15937 414540 16591 414541
rect 15932 413888 15938 414540
rect 16590 413888 16596 414540
rect 15937 413887 16591 413888
rect 19889 412974 20021 412979
rect 19889 412969 19894 412974
rect 20016 412969 20021 412974
rect 19889 412841 20021 412847
rect 576828 411318 576940 417764
rect 578953 417734 579479 417735
rect 578948 417210 578954 417734
rect 579478 417210 579484 417734
rect 578953 417209 579479 417210
rect 578354 414665 578364 414670
rect 578354 414515 578359 414665
rect 578354 414510 578364 414515
rect 578514 414510 578520 414670
rect 576828 411206 581964 411318
rect 582074 411206 584800 411318
rect 20297 410971 20517 410976
rect 19499 410761 20302 410971
rect 20512 410761 20517 410971
rect 19499 409573 19709 410761
rect 20297 410756 20517 410761
rect 583520 410024 584800 410136
rect 13297 409363 19709 409573
rect 13297 394599 13507 409363
rect 582191 409194 582717 409200
rect 582717 408954 582952 409194
rect 582717 408842 584800 408954
rect 582717 408668 582952 408842
rect 582191 408662 582717 408668
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 583520 405296 584800 405408
rect 569970 396573 572430 403252
rect 4463 394389 13507 394599
rect 4463 382107 4673 394389
rect 569965 394115 569971 396573
rect 572429 394115 572435 396573
rect 569970 394114 572430 394115
rect 2385 381976 4673 382107
rect -800 381897 4673 381976
rect -800 381864 2726 381897
rect 2614 381854 2726 381864
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect 9299 371411 9309 371416
rect 9299 371169 9304 371411
rect 9299 371164 9309 371169
rect 9551 371164 9557 371416
rect 10384 365476 36592 390756
rect 52974 370328 52980 374172
rect 56824 370328 56830 374172
rect 13434 346870 13704 365476
rect 13429 346865 13709 346870
rect 13429 346595 13434 346865
rect 13704 346595 13709 346865
rect 13429 346590 13709 346595
rect 11817 345396 11887 345401
rect 13977 345396 14043 345399
rect 11817 345336 11822 345396
rect 11882 345394 14043 345396
rect 11882 345338 13982 345394
rect 14038 345338 14043 345394
rect 11882 345336 14043 345338
rect 11817 345331 11887 345336
rect 13977 345333 14043 345336
rect 18472 343692 18478 343694
rect 15298 343632 18478 343692
rect 14078 343573 14148 343578
rect 14078 343511 14083 343573
rect 14143 343572 14148 343573
rect 15298 343572 15358 343632
rect 18472 343630 18478 343632
rect 18542 343630 18548 343694
rect 14143 343512 15358 343572
rect 14143 343511 14148 343512
rect 14078 343506 14148 343511
rect 16398 341473 17246 341478
rect 16397 341472 17247 341473
rect 14305 341362 14375 341367
rect 14305 341302 14310 341362
rect 14370 341302 14375 341362
rect 14305 341297 14375 341302
rect 14310 340666 14370 341297
rect 14230 340606 14370 340666
rect 16397 340624 16398 341472
rect 17246 340624 17247 341472
rect 16397 340623 17247 340624
rect 16398 340618 17246 340623
rect 9257 340066 9499 340071
rect 9257 339834 9262 340066
rect 9494 339834 9499 340066
rect 9257 339829 9499 339834
rect 14230 339830 14290 340606
rect -800 338710 1870 338754
rect 9262 338710 9494 339829
rect 11442 339702 14314 339830
rect 11442 338710 11570 339702
rect -800 338642 11570 338710
rect 1698 338582 11570 338642
rect 1698 338356 6658 338582
rect 1698 337980 2248 338356
rect 2636 338298 6658 338356
rect 2636 337980 6356 338298
rect 1698 337718 2778 337980
rect -800 337460 480 337572
rect 1698 336765 2074 337718
rect 1693 336391 1699 336765
rect 2073 336391 2079 336765
rect 1698 336390 2074 336391
rect -800 336278 480 336390
rect -800 335096 480 335208
rect 5980 335136 6356 337980
rect 14735 337406 18589 337411
rect 52980 337406 56824 370328
rect 581974 364784 584800 364896
rect 581974 364532 582086 364784
rect 581974 358376 582086 364420
rect 582617 363812 582918 363813
rect 582612 363640 582618 363812
rect 582790 363714 582918 363812
rect 582790 363640 584800 363714
rect 582617 363639 584800 363640
rect 582836 363602 584800 363639
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 583520 358874 584800 358986
rect 581974 358264 583006 358376
rect -800 333914 480 334026
rect 14735 333562 14740 337406
rect 18584 333562 56824 337406
rect 132990 336012 159198 349368
rect 120734 335952 159198 336012
rect 14735 333557 18589 333562
rect -800 332732 480 332844
rect 22866 332378 24484 332383
rect 22866 330770 22871 332378
rect 24479 330770 24484 332378
rect 12106 330691 12238 330696
rect 12106 330686 12111 330691
rect 12233 330686 12238 330691
rect 12106 330570 12238 330576
rect 12239 328544 12517 328549
rect 12239 328276 12244 328544
rect 12512 328276 14670 328544
rect 12239 328271 12517 328276
rect 13410 328222 14670 328276
rect 22866 328222 24484 330770
rect 13410 327704 24484 328222
rect 13452 326611 24484 327704
rect 11768 324843 12628 324849
rect 11768 323988 11773 323993
rect 12623 323988 12628 323993
rect 11768 323983 12628 323988
rect 13452 317662 24356 326611
rect 8337 311290 8439 311295
rect 8336 311289 8440 311290
rect 8336 311187 8337 311289
rect 8439 311187 8440 311289
rect 8336 311186 8440 311187
rect 8337 311181 8439 311186
rect 4887 308208 5487 308213
rect 4887 308203 4892 308208
rect 5482 308203 5487 308208
rect 4887 307607 5487 307613
rect 11703 306480 11913 306485
rect 10638 306280 11708 306480
rect 11908 306280 11913 306480
rect 11703 306275 11913 306280
rect 2721 301936 2731 301941
rect 2721 300636 2726 301936
rect 2721 300631 2731 300636
rect 4031 300631 4037 301941
rect 2857 295534 2959 295539
rect 104 295533 2960 295534
rect 104 295532 2857 295533
rect -800 295431 2857 295532
rect 2959 295431 2960 295533
rect -800 295430 2960 295431
rect -800 295420 480 295430
rect 2857 295425 2959 295430
rect -800 294238 480 294350
rect -800 293056 480 293168
rect 9200 292865 10500 303232
rect 9195 292860 10505 292865
rect -800 291874 480 291986
rect 9195 291560 9200 292860
rect 10500 291560 10505 292860
rect 9195 291555 10505 291560
rect 38176 291680 65700 295542
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 38176 285708 65222 291680
rect 38176 285248 65220 285708
rect 38176 278806 65198 285248
rect 35039 276767 35049 276772
rect 35039 276629 35044 276767
rect 35039 276624 35049 276629
rect 35187 276624 35193 276772
rect 38176 273532 65700 278806
rect 68793 278468 68894 279528
rect 68788 278463 68899 278468
rect 68788 278362 68793 278463
rect 68894 278362 68899 278463
rect 68788 278357 68899 278362
rect 67450 276055 67566 276060
rect 72754 276055 98962 295220
rect 113629 288920 113639 288925
rect 113629 288820 113634 288920
rect 113629 288815 113639 288820
rect 113739 288815 113745 288925
rect 113443 288380 113553 288385
rect 113443 288280 113448 288380
rect 113548 288280 114084 288380
rect 113443 288275 113553 288280
rect 114915 287353 115405 287359
rect 114915 286880 114920 286885
rect 115400 286880 115405 286885
rect 114915 286875 115405 286880
rect 109126 286297 109626 286298
rect 109121 285799 109127 286297
rect 109625 285799 109631 286297
rect 109126 285798 109626 285799
rect 120734 285488 120794 335952
rect 129746 330759 129756 330764
rect 129746 330645 129751 330759
rect 129746 330640 129756 330645
rect 129870 330640 129876 330764
rect 132990 324088 159198 335952
rect 155845 323305 156007 323311
rect 155845 323148 155850 323153
rect 156002 323148 156007 323153
rect 155845 323143 156007 323148
rect 582894 320106 583006 358264
rect 580844 319994 583006 320106
rect 128163 305774 128229 305777
rect 132886 305774 159094 319144
rect 580844 312206 580956 319994
rect 583478 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 582036 313874 582360 313880
rect 582360 313755 583240 313874
rect 583520 313755 584800 313764
rect 582360 313685 584800 313755
rect 582360 313645 583275 313685
rect 583520 313652 584800 313685
rect 582360 313550 583240 313645
rect 582036 313544 582360 313550
rect 580844 312094 583176 312206
rect 128163 305772 159094 305774
rect 128163 305716 128168 305772
rect 128224 305716 159094 305772
rect 128163 305714 159094 305716
rect 128163 305711 128229 305714
rect 131166 299275 131176 299280
rect 131166 299161 131171 299275
rect 131166 299156 131176 299161
rect 131290 299156 131296 299280
rect 132886 293864 159094 305714
rect 204775 307775 219041 307781
rect 199487 293708 199965 293713
rect 199487 293703 199492 293708
rect 199960 293703 199965 293708
rect 582036 300653 582360 300654
rect 582031 300331 582037 300653
rect 582359 300331 582365 300653
rect 582036 300330 582360 300331
rect 579359 295815 579465 295821
rect 579359 295714 579364 295719
rect 579460 295714 579465 295719
rect 579359 295709 579465 295714
rect 581302 295131 581362 296230
rect 581668 295545 581678 295550
rect 581668 295359 581673 295545
rect 581668 295354 581678 295359
rect 581852 295354 581858 295550
rect 581297 295126 581367 295131
rect 581297 295066 581302 295126
rect 581362 295066 581367 295126
rect 581297 295061 581367 295066
rect 583064 293701 583176 312094
rect 583064 293599 583069 293701
rect 583171 293599 583176 293701
rect 583064 293594 583176 293599
rect 204775 293514 204780 293519
rect 219036 293514 219041 293519
rect 204775 293509 219041 293514
rect 199487 293229 199965 293235
rect 581489 290490 581779 290495
rect 581489 290210 581494 290490
rect 581774 290210 581779 290490
rect 581489 290205 581779 290210
rect 107584 285428 120794 285488
rect 107584 283935 107644 285428
rect 110143 285344 110209 285349
rect 110143 285288 110148 285344
rect 110204 285288 110209 285344
rect 110143 285283 110209 285288
rect 110146 285008 110206 285283
rect 111289 285008 111355 285011
rect 110146 285006 111355 285008
rect 110146 284950 111294 285006
rect 111350 284950 111355 285006
rect 110146 284948 111355 284950
rect 111289 284945 111355 284948
rect 111612 284034 111672 284036
rect 113787 284034 113857 284039
rect 111602 283974 113792 284034
rect 113852 283974 113857 284034
rect 107579 283930 107649 283935
rect 107579 283870 107584 283930
rect 107644 283870 107649 283930
rect 107579 283865 107649 283870
rect 109461 283870 109531 283875
rect 111612 283870 111672 283974
rect 113787 283969 113857 283974
rect 109461 283810 109466 283870
rect 109526 283810 111672 283870
rect 109461 283805 109531 283810
rect 110590 278421 110600 278426
rect 110590 278239 110595 278421
rect 110590 278234 110600 278239
rect 110770 278234 110776 278426
rect 110391 277726 110401 277731
rect 110391 277626 110396 277726
rect 110391 277621 110401 277626
rect 110501 277621 110507 277731
rect 67450 275949 67455 276055
rect 67561 275949 98962 276055
rect 67450 275944 67566 275949
rect 68542 273760 68662 273766
rect 68542 273645 68547 273650
rect 68657 273645 68662 273650
rect 68542 273640 68662 273645
rect 38176 273042 65708 273532
rect 66048 273405 66848 273410
rect 66047 273404 66849 273405
rect 6982 258909 33190 269788
rect 38176 269372 65700 273042
rect 66047 272604 66048 273404
rect 66848 272604 66849 273404
rect 66047 272603 66849 272604
rect 66048 272598 66848 272603
rect 72754 269940 98962 275949
rect 133162 275738 159370 290130
rect 577012 289490 577232 289496
rect 577012 289275 577017 289280
rect 577227 289275 577232 289280
rect 577012 289270 577232 289275
rect 580328 289485 580548 289490
rect 580328 289480 580333 289485
rect 580543 289480 580548 289485
rect 580328 289264 580548 289270
rect 581494 288418 581774 290205
rect 573406 288138 581774 288418
rect 573406 287997 573686 288138
rect 573381 287991 573686 287997
rect 573683 287711 573686 287991
rect 573381 287706 573386 287711
rect 573678 287706 573686 287711
rect 573381 287701 573686 287706
rect 573406 287672 573686 287701
rect 581744 287500 582292 287780
rect 217591 287438 217601 287443
rect 199672 282609 200172 284134
rect 199667 282604 200177 282609
rect 199667 282104 199672 282604
rect 200172 282104 200177 282604
rect 199667 282099 200177 282104
rect 217591 279916 217596 287438
rect 217591 279911 217601 279916
rect 225123 279911 225129 287443
rect 108178 275678 159370 275738
rect 107553 274384 107623 274389
rect 108178 274384 108238 275678
rect 107553 274324 107558 274384
rect 107618 274324 108238 274384
rect 109457 274324 109527 274329
rect 107553 274319 107623 274324
rect 109457 274264 109462 274324
rect 109522 274264 127210 274324
rect 109457 274259 109527 274264
rect 104884 269399 104988 269400
rect 40971 268668 41065 268673
rect 41570 268668 41654 269372
rect 104879 269297 104885 269399
rect 104987 269297 104993 269399
rect 104884 269296 104988 269297
rect 119827 269208 120325 269213
rect 119826 269207 120326 269208
rect 119826 268709 119827 269207
rect 120325 268709 120326 269207
rect 119826 268708 120326 268709
rect 119827 268703 120325 268708
rect 40971 268584 40976 268668
rect 41060 268584 41656 268668
rect 87103 268641 87249 268647
rect 83329 268603 83953 268608
rect 69825 268598 83334 268603
rect 40971 268579 41065 268584
rect 69825 267994 69830 268598
rect 70434 267994 83334 268598
rect 69825 267989 83334 267994
rect 83948 267989 83953 268603
rect 87103 268500 87108 268505
rect 87244 268500 87249 268505
rect 87103 268495 87249 268500
rect 110846 268112 111346 268118
rect 83329 267984 83953 267989
rect 68261 267686 82233 267691
rect 68261 267366 68266 267686
rect 68586 267366 82233 267686
rect 68261 267361 82233 267366
rect 69151 266456 69481 267361
rect 70831 267288 70973 267293
rect 70831 267283 70836 267288
rect 70968 267283 70973 267288
rect 70831 267145 70973 267151
rect 36692 264988 36702 264993
rect 36692 264895 36697 264988
rect 36692 264890 36702 264895
rect 36795 264890 36801 264993
rect 43052 262626 46626 263134
rect 37434 260380 37444 260385
rect 37434 260287 37439 260380
rect 37434 260282 37444 260287
rect 37537 260282 37543 260385
rect 33478 258909 33558 258914
rect 6982 258839 33483 258909
rect 33553 258839 33558 258909
rect -800 252398 3586 252510
rect 3698 252398 3704 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect 6982 244508 33190 258839
rect 33478 258834 33558 258839
rect 46118 256656 46626 262626
rect 49859 258900 49869 258905
rect 49859 258744 49864 258900
rect 49859 258739 49869 258744
rect 50025 258739 50031 258905
rect 52064 256656 78272 266456
rect 35443 255778 36087 255783
rect 35443 255144 35448 255778
rect 36082 255144 36087 255778
rect 38630 255277 38734 256294
rect 43204 256148 78272 256656
rect 38630 255183 38635 255277
rect 38729 255183 38734 255277
rect 38630 255178 38734 255183
rect 35443 255139 36087 255144
rect 2726 236473 4026 236474
rect 2721 235175 2727 236473
rect 4025 235175 4031 236473
rect 2726 235174 4026 235175
rect 35448 231397 36082 255139
rect 52064 250438 78272 256148
rect 81903 251329 82233 267361
rect 108424 267612 110846 268112
rect 108424 267275 108924 267612
rect 110846 267606 111346 267612
rect 108424 266785 108429 267275
rect 108919 266785 108924 267275
rect 108424 266208 108924 266785
rect 93350 266037 119558 266208
rect 88654 260959 88982 260964
rect 88653 260958 88983 260959
rect 88653 260630 88654 260958
rect 88982 260630 88983 260958
rect 88653 260629 88983 260630
rect 88654 260624 88982 260629
rect 87441 260510 87511 260515
rect 87441 260440 87446 260510
rect 87506 260505 87511 260510
rect 93350 260505 119564 266037
rect 87506 260445 119564 260505
rect 87506 260440 87511 260445
rect 87441 260435 87511 260440
rect 90579 257328 90897 257333
rect 90579 257020 90584 257328
rect 90892 257020 90897 257328
rect 90579 257015 90897 257020
rect 84749 256528 84923 256529
rect 84744 256356 84750 256528
rect 84922 256356 84928 256528
rect 84749 256355 84923 256356
rect 90584 255997 90892 257015
rect 90584 255699 90589 255997
rect 90887 255699 90892 255997
rect 90584 255694 90892 255699
rect 85334 254618 85340 254802
rect 85514 254797 85524 254802
rect 85519 254623 85524 254797
rect 85514 254618 85524 254623
rect 91664 252561 91674 252566
rect 91664 252443 91669 252561
rect 91664 252438 91674 252443
rect 91792 252438 91798 252566
rect 81093 251307 82233 251329
rect 81093 251197 81153 251307
rect 81275 251197 82233 251307
rect 81093 250999 82233 251197
rect 81093 250438 81423 250999
rect 93350 250438 119564 260445
rect 127150 257334 127210 274264
rect 131600 267887 131610 267892
rect 131600 267773 131605 267887
rect 131600 267768 131610 267773
rect 131724 267768 131730 267892
rect 133162 264850 159370 275678
rect 581644 275247 581922 275252
rect 581644 275145 581649 275247
rect 581751 275145 581922 275247
rect 581644 275140 581922 275145
rect 583488 275140 584800 275252
rect 213025 274928 213035 274933
rect 213025 274817 213030 274928
rect 213025 274812 213035 274817
rect 213146 274812 213152 274933
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 157322 264311 157530 264317
rect 157322 264108 157327 264113
rect 157525 264108 157530 264113
rect 157322 264103 157530 264108
rect 161567 262959 161573 263241
rect 161855 262959 161861 263241
rect 132800 257334 159008 261034
rect 127150 257274 159008 257334
rect 52064 250389 119564 250438
rect 52064 250059 86364 250389
rect 86694 250059 119564 250389
rect 52064 247368 119564 250059
rect 52064 245368 119558 247368
rect 52064 241176 78272 245368
rect 87453 241679 87459 242065
rect 87835 242060 87845 242065
rect 87840 241684 87845 242060
rect 87835 241679 87845 241684
rect 93350 240928 119558 245368
rect 131586 244483 131596 244488
rect 131586 244369 131591 244483
rect 131586 244364 131596 244369
rect 131710 244364 131716 244488
rect 79963 239428 81273 239433
rect 79963 239423 79968 239428
rect 81268 239423 81273 239428
rect 79963 238117 81273 238123
rect 104308 238042 110434 240928
rect 119280 239512 119286 239720
rect 119472 239715 119482 239720
rect 119477 239517 119482 239715
rect 119472 239512 119482 239517
rect 111905 239204 112123 239209
rect 111905 239199 111910 239204
rect 112118 239199 112123 239204
rect 111905 238985 112123 238991
rect 92784 235956 119300 238042
rect 121063 235961 121133 235966
rect 121063 235956 121068 235961
rect 92784 235896 121068 235956
rect 89305 235008 89645 235014
rect 89305 234673 89310 234678
rect 89640 234673 89645 234678
rect 89305 234668 89645 234673
rect 91165 232920 91175 232925
rect 91165 231620 91170 232920
rect 91165 231615 91175 231620
rect 92475 231615 92481 232925
rect 35442 230763 35448 231397
rect 36082 230763 36088 231397
rect 79398 227580 80698 231210
rect 92784 229240 119300 235896
rect 121063 235891 121068 235896
rect 121128 235891 121133 235961
rect 121063 235886 121133 235891
rect 132800 235754 159008 257274
rect 159709 245287 159715 245433
rect 159851 245428 159861 245433
rect 159856 245292 159861 245428
rect 159851 245287 159861 245292
rect 161082 241967 161092 241972
rect 161082 241853 161087 241967
rect 161082 241848 161092 241853
rect 161206 241848 161212 241972
rect 161573 237284 161855 262959
rect 165533 262745 165539 263223
rect 166007 263218 166017 263223
rect 166012 262750 166017 263218
rect 166007 262745 166017 262750
rect 169090 257799 169241 257800
rect 169085 257650 169091 257799
rect 169240 257650 169246 257799
rect 166568 257253 166574 257485
rect 166796 257480 166806 257485
rect 166801 257258 166806 257480
rect 166796 257253 166806 257258
rect 169090 255321 169241 257650
rect 169090 255180 169095 255321
rect 169236 255180 169241 255321
rect 169090 255175 169241 255180
rect 195087 254013 195097 254018
rect 195087 253799 195092 254013
rect 195087 253794 195097 253799
rect 195311 253794 195317 254018
rect 167332 253169 167452 253174
rect 167332 253162 167337 253169
rect 167328 253059 167337 253162
rect 167447 253162 170691 253169
rect 167447 253059 171864 253162
rect 167328 252662 171864 253059
rect 169944 252190 171864 252662
rect 166290 250813 166296 251005
rect 166478 251000 166488 251005
rect 166483 250818 166488 251000
rect 166478 250813 166488 250818
rect 166467 246376 166989 246381
rect 166467 245876 166472 246376
rect 166984 245876 166989 246376
rect 166467 245871 166989 245876
rect 166478 245440 166978 245871
rect 169944 245440 170459 252190
rect 211546 248879 237754 272504
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 582885 269398 583154 269403
rect 582885 269139 582890 269398
rect 583149 269342 583214 269398
rect 583149 269230 584800 269342
rect 583149 269139 583214 269230
rect 582885 269134 583154 269139
rect 166478 245104 170459 245440
rect 163906 245058 170459 245104
rect 163128 244917 170459 245058
rect 210067 248785 237754 248879
rect 163128 243677 170382 244917
rect 163128 243447 163911 243677
rect 164141 243447 170382 243677
rect 163128 242982 170382 243447
rect 161568 237279 161860 237284
rect 161568 236997 161573 237279
rect 161855 236997 161860 237279
rect 161568 236992 161860 236997
rect 92784 228126 119226 229240
rect 124151 228439 124157 228921
rect 124629 228916 124639 228921
rect 124634 228444 124639 228916
rect 124629 228439 124639 228444
rect 84407 227580 85717 227585
rect 92784 227580 119300 228126
rect 5348 227575 84412 227580
rect 5348 226285 5353 227575
rect 6643 226285 84412 227575
rect 5348 226280 84412 226285
rect 85712 226280 119300 227580
rect 84407 226275 85717 226280
rect 92784 225034 119300 226280
rect 139826 225034 141902 225474
rect 163128 225034 165204 242982
rect 179722 225642 182630 225752
rect 179722 225540 187028 225642
rect 187414 225540 188838 225642
rect 179722 225512 188838 225540
rect 181946 225402 188838 225512
rect 186750 225334 187912 225402
rect 186750 225332 187528 225334
rect 92784 224632 172206 225034
rect 92784 224392 177026 224632
rect 92784 223421 176250 224392
rect 92784 223079 168333 223421
rect 168687 223079 176250 223421
rect 92784 222986 176250 223079
rect 92784 222958 172206 222986
rect -800 214888 1660 219688
rect 92784 212868 119300 222958
rect 208912 222170 208922 222175
rect 208912 221956 208917 222170
rect 208912 221951 208922 221956
rect 209136 221951 209142 222175
rect 93018 212742 119226 212868
rect -800 204888 1660 209688
rect 102560 189801 108228 212742
rect 192488 210493 192592 210498
rect 210067 210493 210161 248785
rect 211546 247224 237754 248785
rect 211836 215036 238044 240316
rect 576530 239802 578990 239808
rect 582340 237690 584800 240030
rect 578990 237342 584800 237690
rect 576530 237205 584800 237342
rect 576530 236995 581625 237205
rect 581835 236995 584800 237205
rect 576530 236482 584800 236995
rect 578990 235230 584800 236482
rect 576530 232970 578990 234022
rect 576530 229672 578990 230510
rect 581995 229672 582205 235230
rect 582340 229672 584800 230030
rect 576212 227212 584800 229672
rect 582340 225230 584800 227212
rect 192488 210399 192493 210493
rect 192587 210399 210161 210493
rect 192488 210394 192592 210399
rect 192676 209679 192780 209684
rect 212765 209679 212859 215036
rect 192676 209585 192681 209679
rect 192775 209585 212859 209679
rect 558616 209800 581040 210204
rect 192676 209580 192780 209585
rect 558616 204898 581180 209800
rect 164882 198319 164892 198324
rect 164882 198037 164887 198319
rect 164882 198032 164892 198037
rect 165174 198032 165180 198324
rect 102555 184135 102561 189801
rect 108227 184135 108233 189801
rect 102560 184134 108228 184135
rect 582340 194750 584800 196230
rect 581180 192290 584800 194750
rect 582340 191430 584800 192290
rect 582340 184750 584800 186230
rect 581180 182334 584800 184750
rect 558616 182328 584800 182334
rect 578720 182290 584800 182328
rect 582340 181430 584800 182290
rect -800 172888 1660 177688
rect -800 162888 1660 167688
rect 582340 146830 584800 151630
rect 582340 136830 584800 141630
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 480 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< rmetal3 >>
rect 583234 589452 583356 589596
rect 12902 462398 13008 462510
rect 581964 411202 582074 411328
rect 581974 364420 582086 364532
<< via3 >>
rect 583004 589472 583116 589584
rect 568898 497457 569048 497462
rect 568898 497307 568903 497457
rect 568903 497307 569048 497457
rect 568898 497302 569048 497307
rect 576659 496070 576903 496075
rect 576659 495826 576898 496070
rect 576898 495826 576903 496070
rect 576659 495821 576903 495826
rect 579365 483287 581823 485745
rect 18616 462398 18728 462510
rect 579365 445635 581823 448093
rect 15187 431528 15767 431533
rect 15187 430948 15762 431528
rect 15762 430948 15767 431528
rect 15187 430943 15767 430948
rect 576267 424394 576367 424399
rect 576267 424294 576272 424394
rect 576272 424294 576367 424394
rect 576267 424289 576367 424294
rect 578927 422614 579102 422619
rect 578927 422439 579097 422614
rect 579097 422439 579102 422614
rect 578927 422434 579102 422439
rect 27814 417016 28662 417020
rect 27814 416176 27818 417016
rect 27818 416176 28658 417016
rect 28658 416176 28662 417016
rect 27814 416172 28662 416176
rect 572817 416270 573027 416275
rect 572817 416075 572822 416270
rect 572822 416075 573022 416270
rect 573022 416075 573027 416270
rect 15938 414536 16590 414540
rect 15938 413892 15942 414536
rect 15942 413892 16586 414536
rect 16586 413892 16590 414536
rect 15938 413888 16590 413892
rect 19889 412852 19894 412969
rect 19894 412852 20016 412969
rect 20016 412852 20021 412969
rect 19889 412847 20021 412852
rect 578954 417730 579478 417734
rect 578954 417214 578958 417730
rect 578958 417214 579474 417730
rect 579474 417214 579478 417730
rect 578954 417210 579478 417214
rect 578364 414665 578514 414670
rect 578364 414515 578509 414665
rect 578509 414515 578514 414665
rect 578364 414510 578514 414515
rect 582191 408668 582717 409194
rect 569971 394115 572429 396573
rect 9309 371411 9551 371416
rect 9309 371169 9546 371411
rect 9546 371169 9551 371411
rect 9309 371164 9551 371169
rect 52980 370328 56824 374172
rect 18478 343630 18542 343694
rect 16398 341468 17246 341472
rect 16398 340628 16402 341468
rect 16402 340628 17242 341468
rect 17242 340628 17246 341468
rect 16398 340624 17246 340628
rect 1699 336391 2073 336765
rect 582618 363640 582790 363812
rect 12106 330581 12111 330686
rect 12111 330581 12233 330686
rect 12233 330581 12238 330686
rect 12106 330576 12238 330581
rect 11768 324838 12628 324843
rect 11768 323993 11773 324838
rect 11773 323993 12623 324838
rect 12623 323993 12628 324838
rect 8337 311285 8439 311289
rect 8337 311191 8341 311285
rect 8341 311191 8435 311285
rect 8435 311191 8439 311285
rect 8337 311187 8439 311191
rect 4887 307618 4892 308203
rect 4892 307618 5482 308203
rect 5482 307618 5487 308203
rect 4887 307613 5487 307618
rect 2731 301936 4031 301941
rect 2731 300636 4026 301936
rect 4026 300636 4031 301936
rect 2731 300631 4031 300636
rect 2857 295431 2959 295533
rect 35049 276767 35187 276772
rect 35049 276629 35182 276767
rect 35182 276629 35187 276767
rect 35049 276624 35187 276629
rect 113639 288920 113739 288925
rect 113639 288820 113734 288920
rect 113734 288820 113739 288920
rect 113639 288815 113739 288820
rect 114915 287348 115405 287353
rect 114915 286885 114920 287348
rect 114920 286885 115400 287348
rect 115400 286885 115405 287348
rect 109127 286293 109625 286297
rect 109127 285803 109131 286293
rect 109131 285803 109621 286293
rect 109621 285803 109625 286293
rect 109127 285799 109625 285803
rect 129756 330759 129870 330764
rect 129756 330645 129865 330759
rect 129865 330645 129870 330759
rect 129756 330640 129870 330645
rect 155845 323300 156007 323305
rect 155845 323153 155850 323300
rect 155850 323153 156002 323300
rect 156002 323153 156007 323300
rect 582036 313550 582360 313874
rect 131176 299275 131290 299280
rect 131176 299161 131285 299275
rect 131285 299161 131290 299275
rect 131176 299156 131290 299161
rect 204775 307770 219041 307775
rect 199487 293240 199492 293703
rect 199492 293240 199960 293703
rect 199960 293240 199965 293703
rect 204775 293519 204780 307770
rect 204780 293519 219036 307770
rect 219036 293519 219041 307770
rect 582037 300649 582359 300653
rect 582037 300335 582041 300649
rect 582041 300335 582355 300649
rect 582355 300335 582359 300649
rect 582037 300331 582359 300335
rect 579359 295810 579465 295815
rect 579359 295719 579364 295810
rect 579364 295719 579460 295810
rect 579460 295719 579465 295810
rect 581678 295545 581852 295550
rect 581678 295359 581847 295545
rect 581847 295359 581852 295545
rect 581678 295354 581852 295359
rect 199487 293235 199965 293240
rect 110600 278421 110770 278426
rect 110600 278239 110765 278421
rect 110765 278239 110770 278421
rect 110600 278234 110770 278239
rect 110401 277726 110501 277731
rect 110401 277626 110496 277726
rect 110496 277626 110501 277726
rect 110401 277621 110501 277626
rect 68542 273755 68662 273760
rect 68542 273650 68547 273755
rect 68547 273650 68657 273755
rect 68657 273650 68662 273755
rect 66048 273400 66848 273404
rect 66048 272608 66052 273400
rect 66052 272608 66844 273400
rect 66844 272608 66848 273400
rect 66048 272604 66848 272608
rect 577012 289485 577232 289490
rect 577012 289280 577017 289485
rect 577017 289280 577227 289485
rect 577227 289280 577232 289485
rect 580328 289275 580333 289480
rect 580333 289275 580543 289480
rect 580543 289275 580548 289480
rect 580328 289270 580548 289275
rect 573381 287986 573683 287991
rect 573381 287711 573386 287986
rect 573386 287711 573678 287986
rect 573678 287711 573683 287986
rect 217601 287438 225123 287443
rect 217601 279916 225118 287438
rect 225118 279916 225123 287438
rect 217601 279911 225123 279916
rect 104885 269395 104987 269399
rect 104885 269301 104889 269395
rect 104889 269301 104983 269395
rect 104983 269301 104987 269395
rect 104885 269297 104987 269301
rect 119827 269203 120325 269207
rect 119827 268713 119831 269203
rect 119831 268713 120321 269203
rect 120321 268713 120325 269203
rect 119827 268709 120325 268713
rect 87103 268636 87249 268641
rect 87103 268505 87108 268636
rect 87108 268505 87244 268636
rect 87244 268505 87249 268636
rect 70831 267156 70836 267283
rect 70836 267156 70968 267283
rect 70968 267156 70973 267283
rect 70831 267151 70973 267156
rect 36702 264988 36795 264993
rect 36702 264895 36790 264988
rect 36790 264895 36795 264988
rect 36702 264890 36795 264895
rect 37444 260380 37537 260385
rect 37444 260287 37532 260380
rect 37532 260287 37537 260380
rect 37444 260282 37537 260287
rect 3586 252398 3698 252510
rect 49869 258900 50025 258905
rect 49869 258744 50020 258900
rect 50020 258744 50025 258900
rect 49869 258739 50025 258744
rect 2727 236469 4025 236473
rect 2727 235179 2731 236469
rect 2731 235179 4021 236469
rect 4021 235179 4025 236469
rect 2727 235175 4025 235179
rect 110846 267612 111346 268112
rect 88654 260954 88982 260958
rect 88654 260634 88658 260954
rect 88658 260634 88978 260954
rect 88978 260634 88982 260954
rect 88654 260630 88982 260634
rect 84750 256524 84922 256528
rect 84750 256360 84754 256524
rect 84754 256360 84918 256524
rect 84918 256360 84922 256524
rect 84750 256356 84922 256360
rect 85340 254797 85514 254802
rect 85340 254623 85345 254797
rect 85345 254623 85514 254797
rect 85340 254618 85514 254623
rect 91674 252561 91792 252566
rect 91674 252443 91787 252561
rect 91787 252443 91792 252561
rect 91674 252438 91792 252443
rect 131610 267887 131724 267892
rect 131610 267773 131719 267887
rect 131719 267773 131724 267887
rect 131610 267768 131724 267773
rect 213035 274928 213146 274933
rect 213035 274817 213141 274928
rect 213141 274817 213146 274928
rect 213035 274812 213146 274817
rect 157322 264306 157530 264311
rect 157322 264113 157327 264306
rect 157327 264113 157525 264306
rect 157525 264113 157530 264306
rect 161573 262959 161855 263241
rect 87459 242060 87835 242065
rect 87459 241684 87464 242060
rect 87464 241684 87835 242060
rect 87459 241679 87835 241684
rect 131596 244483 131710 244488
rect 131596 244369 131705 244483
rect 131705 244369 131710 244483
rect 131596 244364 131710 244369
rect 79963 238128 79968 239423
rect 79968 238128 81268 239423
rect 81268 238128 81273 239423
rect 79963 238123 81273 238128
rect 119286 239715 119472 239720
rect 119286 239517 119291 239715
rect 119291 239517 119472 239715
rect 119286 239512 119472 239517
rect 111905 238996 111910 239199
rect 111910 238996 112118 239199
rect 112118 238996 112123 239199
rect 111905 238991 112123 238996
rect 89305 235003 89645 235008
rect 89305 234678 89310 235003
rect 89310 234678 89640 235003
rect 89640 234678 89645 235003
rect 91175 232920 92475 232925
rect 91175 231620 92470 232920
rect 92470 231620 92475 232920
rect 91175 231615 92475 231620
rect 35448 230763 36082 231397
rect 159715 245428 159851 245433
rect 159715 245292 159720 245428
rect 159720 245292 159851 245428
rect 159715 245287 159851 245292
rect 161092 241967 161206 241972
rect 161092 241853 161201 241967
rect 161201 241853 161206 241967
rect 161092 241848 161206 241853
rect 165539 263218 166007 263223
rect 165539 262750 165544 263218
rect 165544 262750 166007 263218
rect 165539 262745 166007 262750
rect 169091 257650 169240 257799
rect 166574 257480 166796 257485
rect 166574 257258 166579 257480
rect 166579 257258 166796 257480
rect 166574 257253 166796 257258
rect 195097 254013 195311 254018
rect 195097 253799 195306 254013
rect 195306 253799 195311 254013
rect 195097 253794 195311 253799
rect 166296 251000 166478 251005
rect 166296 250818 166301 251000
rect 166301 250818 166478 251000
rect 166296 250813 166478 250818
rect 124157 228916 124629 228921
rect 124157 228444 124162 228916
rect 124162 228444 124629 228916
rect 124157 228439 124629 228444
rect 208922 222170 209136 222175
rect 208922 221956 209131 222170
rect 209131 221956 209136 222170
rect 208922 221951 209136 221956
rect 576530 237342 578990 239802
rect 576530 234022 578990 236482
rect 576530 230510 578990 232970
rect 164892 198319 165174 198324
rect 164892 198037 165169 198319
rect 165169 198037 165174 198319
rect 164892 198032 165174 198037
rect 102561 184135 108227 189801
rect 558616 182334 581180 204898
<< metal4 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 583003 589584 583117 589585
rect 583003 589472 583004 589584
rect 583116 589472 583117 589584
rect 583003 589471 583117 589472
rect 583004 557546 583116 589471
rect 579176 557434 583116 557546
rect 566028 497457 567908 502966
rect 579176 500162 579288 557434
rect 579176 500050 580656 500162
rect 568897 497462 569049 497463
rect 568897 497457 568898 497462
rect 566028 497307 568898 497457
rect 566028 492660 567908 497307
rect 568897 497302 568898 497307
rect 569048 497302 569049 497462
rect 568897 497301 569049 497302
rect 568630 492660 575292 492690
rect 566028 490230 575292 492660
rect 18615 462510 18729 462511
rect 18615 462398 18616 462510
rect 18728 462398 18729 462510
rect 18615 462397 18729 462398
rect 18616 458049 18728 462397
rect 16561 435114 70222 458049
rect 17064 432382 22670 435114
rect 15186 431533 15768 431534
rect 15186 430943 15187 431533
rect 15767 431528 15768 431533
rect 15767 430948 18104 431528
rect 15767 430943 15768 430948
rect 15186 430942 15768 430943
rect 27813 417020 28663 417021
rect 27813 416172 27814 417020
rect 28662 416172 28663 417020
rect 27813 416171 28663 416172
rect 2969 414540 16591 414541
rect 2969 413888 15938 414540
rect 16590 413888 16591 414540
rect 2969 413887 16591 413888
rect 1698 336765 2074 336766
rect 1698 336391 1699 336765
rect 2073 336391 2074 336765
rect 1698 336390 2074 336391
rect 2969 308161 3623 413887
rect 19888 412969 20022 412970
rect 19888 412847 19889 412969
rect 20021 412847 20022 412969
rect 19888 412846 20022 412847
rect 19894 411255 20016 412846
rect 19677 409489 20103 411255
rect 19677 409063 20356 409489
rect 5811 350143 6661 401641
rect 19930 390434 20356 409063
rect 47287 397107 70222 435114
rect 572832 424394 575292 490230
rect 579364 485745 581824 485746
rect 579364 483287 579365 485745
rect 581823 483287 581824 485745
rect 579364 483286 581824 483287
rect 579364 448093 581824 448094
rect 579364 445635 579365 448093
rect 581823 445635 581824 448093
rect 579364 445634 581824 445635
rect 576266 424399 576368 424400
rect 576266 424394 576267 424399
rect 572832 424294 576267 424394
rect 572832 419396 575292 424294
rect 576266 424289 576267 424294
rect 576367 424289 576368 424399
rect 576266 424288 576368 424289
rect 570144 416936 575292 419396
rect 578953 417734 582717 417735
rect 578953 417210 578954 417734
rect 579478 417210 582717 417734
rect 578953 417209 582717 417210
rect 570144 416275 572604 416936
rect 572816 416275 573028 416276
rect 570144 416075 572817 416275
rect 573027 416075 573028 416275
rect 570144 410072 572604 416075
rect 572816 416074 573028 416075
rect 570144 407612 577630 410072
rect 582191 409195 582717 417209
rect 582190 409194 582718 409195
rect 582190 408668 582191 409194
rect 582717 408668 582718 409194
rect 582190 408667 582718 408668
rect 47287 374172 287119 397107
rect 569970 396573 572430 396574
rect 569970 394115 569971 396573
rect 572429 394115 572430 396573
rect 569970 394114 572430 394115
rect 9308 371416 9552 371417
rect 9308 371164 9309 371416
rect 9551 371411 9552 371416
rect 9656 371411 11701 371449
rect 9551 371207 11701 371411
rect 9551 371169 9905 371207
rect 9551 371164 9552 371169
rect 9308 371163 9552 371164
rect 47287 370328 52980 374172
rect 56824 370328 287119 374172
rect 47287 369733 287119 370328
rect 13296 364278 14220 366462
rect 19350 364278 20274 368248
rect 26142 364278 27066 366774
rect 33732 364278 34656 366950
rect 13296 363354 34656 364278
rect 29434 359906 184808 361046
rect 5811 349293 10857 350143
rect 10007 339165 10857 349293
rect 29434 343808 30574 359906
rect 135744 350213 156215 350659
rect 135744 349008 136190 350213
rect 142571 348937 143017 350213
rect 149061 348363 149507 350213
rect 155769 348887 156215 350213
rect 18477 343694 18543 343695
rect 18477 343630 18478 343694
rect 18542 343692 18543 343694
rect 20456 343692 30574 343808
rect 18542 343632 30574 343692
rect 18542 343630 18543 343632
rect 18477 343629 18543 343630
rect 20456 342668 30574 343632
rect 16397 341472 17247 341473
rect 16397 340624 16398 341472
rect 17246 340624 17247 341472
rect 16397 339165 17247 340624
rect 10007 338315 17247 339165
rect 8357 330253 9207 331641
rect 11773 330686 12623 338315
rect 11773 330576 12106 330686
rect 12238 330576 12623 330686
rect 129755 330764 129871 330765
rect 129755 330640 129756 330764
rect 129870 330759 129871 330764
rect 136101 330759 136215 331905
rect 129870 330645 136215 330759
rect 129870 330640 129871 330645
rect 129755 330639 129871 330640
rect 11773 330253 12623 330576
rect 8357 329403 12623 330253
rect 11773 324844 12623 329403
rect 183668 327650 184808 359906
rect 183668 326510 247292 327650
rect 11767 324843 12629 324844
rect 11767 323993 11768 324843
rect 12628 323993 12629 324843
rect 11767 323992 12629 323993
rect 155850 323306 156002 324558
rect 155844 323305 156008 323306
rect 155844 323153 155845 323305
rect 156007 323153 156008 323305
rect 155844 323152 156008 323153
rect 135754 319583 156153 319945
rect 135754 318804 136116 319583
rect 142435 318691 142797 319583
rect 148981 318307 149343 319583
rect 155791 318869 156153 319583
rect 15920 316928 16024 317774
rect 21542 316928 21646 317992
rect 12382 316824 21646 316928
rect 12382 311290 12486 316824
rect 8336 311289 12486 311290
rect 8336 311187 8337 311289
rect 8439 311187 12486 311289
rect 8336 311186 12486 311187
rect 4886 308203 5488 308204
rect 4093 308161 4887 308203
rect 2969 307613 4887 308161
rect 5487 307613 5488 308203
rect 2969 307507 4715 307613
rect 4886 307612 5488 307613
rect 4093 306393 4683 307507
rect 4093 305803 5913 306393
rect 2730 301941 4032 301942
rect 2730 300631 2731 301941
rect 4031 301936 4032 301941
rect 4031 300636 6946 301936
rect 4031 300631 4032 300636
rect 2730 300630 4032 300631
rect 12382 295534 12486 311186
rect 131175 299280 131291 299281
rect 131175 299156 131176 299280
rect 131290 299275 131291 299280
rect 131290 299161 133753 299275
rect 131290 299156 131291 299161
rect 131175 299155 131291 299156
rect 2856 295533 12486 295534
rect 2856 295431 2857 295533
rect 2959 295431 12486 295533
rect 2856 295430 12486 295431
rect 75530 296307 96255 297037
rect 75530 294300 76260 296307
rect 82057 294017 82787 296307
rect 88677 294539 89407 296307
rect 95525 294163 96255 296307
rect 157235 291660 157386 294379
rect 199486 293703 199966 293704
rect 199486 293235 199487 293703
rect 199965 293235 199966 293703
rect 204774 293519 204775 293520
rect 219041 293519 219042 293520
rect 204774 293518 219042 293519
rect 199486 293234 199966 293235
rect 157235 291509 169241 291660
rect 136028 290593 156431 290999
rect 136028 289862 136434 290593
rect 142533 289337 142939 290593
rect 149169 289659 149575 290593
rect 156025 289807 156431 290593
rect 113638 288925 113740 288926
rect 113638 288815 113639 288925
rect 113739 288920 113740 288925
rect 113739 288820 114340 288920
rect 113739 288815 113740 288820
rect 113638 288814 113740 288815
rect 114926 287354 115394 288968
rect 114914 287353 115406 287354
rect 114914 286885 114915 287353
rect 115405 287346 115406 287353
rect 121232 287346 122842 287361
rect 115405 286885 122842 287346
rect 114914 286884 122842 286885
rect 114926 286878 122842 286884
rect 109126 286297 109626 286298
rect 109126 285799 109127 286297
rect 109625 285799 109626 286297
rect 109126 285798 109626 285799
rect 121232 285823 122842 286878
rect 35048 276772 35188 276773
rect 35048 276624 35049 276772
rect 35187 276767 35188 276772
rect 35187 276629 39249 276767
rect 35187 276624 35188 276629
rect 35048 276623 35188 276624
rect 68547 273761 68657 280113
rect 68541 273760 68663 273761
rect 68541 273650 68542 273760
rect 68662 273650 68663 273760
rect 68541 273649 68663 273650
rect 66047 273404 66849 273405
rect 64136 273264 64786 273324
rect 66047 272604 66048 273404
rect 66848 272604 66849 273404
rect 41930 269055 42732 270580
rect 48071 269055 48873 270489
rect 54809 269055 55611 270559
rect 61505 269055 62307 270475
rect 66047 269055 66849 272604
rect 41930 268253 66849 269055
rect 87108 268642 87244 270510
rect 95578 269400 95682 270056
rect 95578 269399 104988 269400
rect 95578 269297 104885 269399
rect 104987 269297 104988 269399
rect 95578 269296 104988 269297
rect 119826 269207 120326 269208
rect 119826 268709 119827 269207
rect 120325 268709 120326 269207
rect 119826 268708 120326 268709
rect 87102 268641 87250 268642
rect 87102 268505 87103 268641
rect 87249 268505 87250 268641
rect 87102 268504 87250 268505
rect 110845 267612 110846 267613
rect 111346 267612 111347 267613
rect 110845 267611 111347 267612
rect 70830 267283 70974 267284
rect 70830 267151 70831 267283
rect 70973 267151 70974 267283
rect 70830 267150 70974 267151
rect 70836 266777 70968 267150
rect 121232 266868 122842 284213
rect 131609 267892 131725 267893
rect 131609 267768 131610 267892
rect 131724 267887 131725 267892
rect 131724 267773 134495 267887
rect 131724 267768 131725 267773
rect 131609 267767 131725 267768
rect 56285 266603 80483 266777
rect 56285 265329 56459 266603
rect 61887 265593 62061 266603
rect 68223 265957 68397 266603
rect 74833 265947 75007 266603
rect 76587 265633 76761 266603
rect 36701 264993 36796 264994
rect 36701 264890 36702 264993
rect 36795 264988 36796 264993
rect 36795 264895 38534 264988
rect 36795 264890 36796 264895
rect 36701 264889 36796 264890
rect 37443 260385 37538 260386
rect 37443 260282 37444 260385
rect 37537 260380 37538 260385
rect 37537 260287 38304 260380
rect 37537 260282 37538 260287
rect 37443 260281 37538 260282
rect 49868 258905 50026 258906
rect 49868 258739 49869 258905
rect 50025 258900 50026 258905
rect 50025 258744 52928 258900
rect 50025 258739 50026 258744
rect 49868 258738 50026 258739
rect 3585 252510 3699 252511
rect 3585 252398 3586 252510
rect 3698 252398 7316 252510
rect 3585 252397 3699 252398
rect 8050 242795 10232 246068
rect 15731 242795 17913 247381
rect 22231 242795 24413 248005
rect 29309 242795 31491 248137
rect 8050 240613 31491 242795
rect 40718 237144 42018 257634
rect 80309 254797 80483 266603
rect 121232 266400 128674 266868
rect 121232 263400 122842 266400
rect 157327 264312 157525 265319
rect 157321 264311 157531 264312
rect 157321 264113 157322 264311
rect 157530 264113 157531 264311
rect 157321 264112 157531 264113
rect 121232 262970 128992 263400
rect 121298 262932 128992 262970
rect 129460 263241 165326 263400
rect 129460 262959 161573 263241
rect 161855 263218 165326 263241
rect 165538 263223 166008 263224
rect 165538 263218 165539 263223
rect 161855 262959 165539 263218
rect 129460 262932 165539 262959
rect 164858 262750 165539 262932
rect 164858 262178 165376 262750
rect 165538 262745 165539 262750
rect 166007 262745 166008 263223
rect 165538 262744 166008 262745
rect 135616 261546 155798 261910
rect 88653 260958 88983 260959
rect 88653 260630 88654 260958
rect 88982 260630 88983 260958
rect 135616 260654 135980 261546
rect 88653 260629 88983 260630
rect 142224 260560 142588 261546
rect 148858 260542 149222 261546
rect 155434 260674 155798 261546
rect 164908 257480 165376 262178
rect 169090 257799 169241 291509
rect 199492 287746 199960 293234
rect 217600 287443 217602 287444
rect 217600 279911 217601 287443
rect 217600 279910 217602 279911
rect 214542 275162 215682 275264
rect 213034 274933 213147 274934
rect 213034 274812 213035 274933
rect 213146 274928 213147 274933
rect 214542 274928 234842 275162
rect 213146 274817 234842 274928
rect 213146 274812 213147 274817
rect 213034 274811 213147 274812
rect 214542 274022 234842 274817
rect 214542 270806 215682 274022
rect 220694 270922 221834 274022
rect 227710 270982 228850 274022
rect 233702 271068 234842 274022
rect 169090 257650 169091 257799
rect 169240 257650 169241 257799
rect 169090 257649 169241 257650
rect 166573 257485 166797 257486
rect 166573 257480 166574 257485
rect 164908 257258 166574 257480
rect 84850 256529 84910 256532
rect 84749 256528 84923 256529
rect 84749 256356 84750 256528
rect 84922 256356 84923 256528
rect 84749 254797 84923 256356
rect 85339 254802 85515 254803
rect 85339 254797 85340 254802
rect 80309 254623 85340 254797
rect 85339 254618 85340 254623
rect 85514 254618 85515 254802
rect 85339 254617 85515 254618
rect 91673 252566 91793 252567
rect 91673 252438 91674 252566
rect 91792 252561 91793 252566
rect 91792 252443 93773 252561
rect 91792 252438 91793 252443
rect 91673 252437 91793 252438
rect 164908 251000 165376 257258
rect 166324 257253 166574 257258
rect 166796 257338 166797 257485
rect 166796 257314 168828 257338
rect 166796 257253 170244 257314
rect 166324 257238 170244 257253
rect 168796 257214 170244 257238
rect 170144 256848 170244 257214
rect 170144 256748 171720 256848
rect 195096 254018 195312 254019
rect 195096 253794 195097 254018
rect 195311 254013 195312 254018
rect 195311 253799 216095 254013
rect 195311 253794 195312 253799
rect 195096 253793 195312 253794
rect 166295 251005 166479 251006
rect 166295 251000 166296 251005
rect 164908 250818 166296 251000
rect 164908 250686 165376 250818
rect 166295 250813 166296 250818
rect 166478 250813 166479 251005
rect 166295 250812 166479 250813
rect 159714 245433 159852 245434
rect 159714 245287 159715 245433
rect 159851 245287 159852 245433
rect 159714 245286 159852 245287
rect 131595 244488 131711 244489
rect 131595 244364 131596 244488
rect 131710 244483 131711 244488
rect 131710 244369 134153 244483
rect 131710 244364 131711 244369
rect 131595 244363 131711 244364
rect 96338 240376 96442 241032
rect 102920 240376 103024 241630
rect 109586 240376 109690 241630
rect 116232 240376 116336 241214
rect 96338 240272 116336 240376
rect 118441 239709 118627 241249
rect 119285 239720 119473 239721
rect 119285 239709 119286 239720
rect 118441 239523 119286 239709
rect 119285 239512 119286 239523
rect 119472 239512 119473 239720
rect 119285 239511 119473 239512
rect 79962 239423 81274 239424
rect 79962 238123 79963 239423
rect 81273 238123 81274 239423
rect 111904 239199 112124 239200
rect 111904 238991 111905 239199
rect 112123 238991 112124 239199
rect 111904 238990 112124 238991
rect 79962 238122 81274 238123
rect 2276 237062 79734 237144
rect 79968 237062 81268 238122
rect 111910 237646 112118 238990
rect 2276 236473 81268 237062
rect 2276 235175 2727 236473
rect 4025 235762 81268 236473
rect 4025 235175 79896 235762
rect 2276 232472 79896 235175
rect 156574 235114 156710 236780
rect 159715 235114 159851 245286
rect 246152 242144 247292 326510
rect 161091 241972 161207 241973
rect 161091 241848 161092 241972
rect 161206 241967 161207 241972
rect 161206 241853 165849 241967
rect 161206 241848 161207 241853
rect 161091 241847 161207 241848
rect 214658 241004 247292 242144
rect 259745 322855 287119 369733
rect 259745 258024 287119 295481
rect 575170 289490 577630 407612
rect 582617 363812 582791 363813
rect 582617 363640 582618 363812
rect 582790 363640 582791 363812
rect 582035 313874 582361 313875
rect 582035 313550 582036 313874
rect 582360 313550 582361 313874
rect 582035 313549 582361 313550
rect 582036 300653 582360 313549
rect 582036 300331 582037 300653
rect 582359 300331 582360 300653
rect 582036 300330 582360 300331
rect 579364 295816 579460 296378
rect 579358 295815 579466 295816
rect 579358 295719 579359 295815
rect 579465 295719 579466 295815
rect 579358 295718 579466 295719
rect 581677 295550 581853 295551
rect 581677 295354 581678 295550
rect 581852 295539 581853 295550
rect 582617 295539 582791 363640
rect 581852 295365 582791 295539
rect 581852 295354 581853 295365
rect 581677 295353 581853 295354
rect 575170 289280 577012 289490
rect 577232 289280 577630 289490
rect 575170 288290 577630 289280
rect 580327 289480 580549 289481
rect 580327 289270 580328 289480
rect 580548 289270 580549 289480
rect 580327 289269 580549 289270
rect 575170 285830 578990 288290
rect 580333 287881 580543 289269
rect 576530 258024 578990 285830
rect 214658 238652 215798 241004
rect 220548 239500 221688 241004
rect 227388 238564 228528 241004
rect 233776 238534 234916 241004
rect 259745 239802 579141 258024
rect 156574 234978 159851 235114
rect 259745 237342 576530 239802
rect 578990 237342 579141 239802
rect 259745 236482 579141 237342
rect 89304 234678 89305 234679
rect 89645 234678 89646 234679
rect 89304 234677 89646 234678
rect 259745 234022 576530 236482
rect 578990 234022 579141 236482
rect 259745 232970 579141 234022
rect 91174 232925 92476 232926
rect 2276 232004 79734 232472
rect 35447 231397 35449 231398
rect 35447 230763 35448 231397
rect 35447 230762 35449 230763
rect 74594 199240 79734 232004
rect 91174 231615 91175 232925
rect 92475 232920 92476 232925
rect 92475 231620 94520 232920
rect 92475 231615 92476 231620
rect 91174 231614 92476 231615
rect 93220 212356 94520 231620
rect 259745 230650 576530 232970
rect 124156 228921 124630 228922
rect 124156 228916 124157 228921
rect 119944 228444 124157 228916
rect 102234 212356 103534 214586
rect 108308 212356 109608 214794
rect 115456 212518 116756 215042
rect 120048 212518 120520 228444
rect 124156 228439 124157 228444
rect 124629 228439 124630 228921
rect 124156 228438 124630 228439
rect 208921 222175 209137 222176
rect 208921 221951 208922 222175
rect 209136 222170 209137 222175
rect 209136 221956 213001 222170
rect 209136 221951 209137 221956
rect 208921 221950 209137 221951
rect 115456 212356 120520 212518
rect 93220 212046 120520 212356
rect 93220 211056 116756 212046
rect 259745 204323 287119 230650
rect 569978 230510 576530 230650
rect 578990 230650 579141 232970
rect 578990 230510 578991 230650
rect 576529 230509 578991 230510
rect 126745 199240 287119 204323
rect 74594 194100 129060 199240
rect 134200 198324 287119 199240
rect 134200 198032 164892 198324
rect 165174 198032 287119 198324
rect 134200 194100 287119 198032
rect 102560 189801 108228 189802
rect 102560 184135 102561 189801
rect 108227 184135 108228 189801
rect 102560 184134 108228 184135
rect 126745 176949 287119 194100
rect 558615 182334 558616 182335
rect 581180 182334 581181 182335
rect 558615 182333 581181 182334
rect 259745 175507 287119 176949
<< via4 >>
rect 580656 499946 580976 500266
rect 576621 496075 576941 496108
rect 576621 495821 576659 496075
rect 576659 495821 576903 496075
rect 576903 495821 576941 496075
rect 576621 495788 576941 495821
rect 27837 416195 28639 416997
rect 1722 336414 2050 336742
rect 5811 401641 6661 402491
rect 579388 483310 581800 485722
rect 579388 445658 581800 448070
rect 578855 422619 579175 422687
rect 578855 422434 578927 422619
rect 578927 422434 579102 422619
rect 579102 422434 579175 422619
rect 578855 422367 579175 422434
rect 578279 414670 578599 414750
rect 578279 414510 578364 414670
rect 578364 414510 578514 414670
rect 578514 414510 578599 414670
rect 578279 414430 578599 414510
rect 569994 394138 572406 396550
rect 204774 307775 219042 307776
rect 204774 293520 204775 307775
rect 204775 293520 219041 307775
rect 219041 293520 219042 307775
rect 109150 285822 109602 286274
rect 121232 284213 122842 285823
rect 110525 278426 110845 278490
rect 110525 278234 110600 278426
rect 110600 278234 110770 278426
rect 110770 278234 110845 278426
rect 110525 278170 110845 278234
rect 110291 277731 110611 277836
rect 110291 277621 110401 277731
rect 110401 277621 110501 277731
rect 110501 277621 110611 277731
rect 110291 277516 110611 277621
rect 119850 268732 120302 269184
rect 110845 268112 111347 268113
rect 110845 267613 110846 268112
rect 110846 267613 111346 268112
rect 111346 267613 111347 268112
rect 128674 266400 129142 266868
rect 128992 262932 129460 263400
rect 88677 260653 88959 260935
rect 217602 287443 225124 287444
rect 217602 279911 225123 287443
rect 225123 279911 225124 287443
rect 217602 279910 225124 279911
rect 87458 242065 87836 242066
rect 87458 241679 87459 242065
rect 87459 241679 87835 242065
rect 87835 241679 87836 242065
rect 87458 241678 87836 241679
rect 259745 295481 287119 322855
rect 573372 287991 573692 288011
rect 573372 287711 573381 287991
rect 573381 287711 573683 287991
rect 573683 287711 573692 287991
rect 573372 287691 573692 287711
rect 89304 235008 89646 235009
rect 89304 234679 89305 235008
rect 89305 234679 89645 235008
rect 89645 234679 89646 235008
rect 35449 231397 36083 231398
rect 35449 230763 36082 231397
rect 36082 230763 36083 231397
rect 35449 230762 36083 230763
rect 129060 194100 134200 199240
rect 102584 184158 108204 189778
rect 558615 204898 581181 204899
rect 558615 182335 558616 204898
rect 558616 182335 581180 204898
rect 581180 182335 581181 204898
<< metal5 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 580632 500266 581000 500290
rect 580632 499946 580656 500266
rect 580976 499946 581000 500266
rect 580632 499922 581000 499946
rect 580656 498444 580976 499922
rect 576597 496108 576965 496132
rect 579364 496108 581824 498444
rect 576597 495788 576621 496108
rect 576941 495788 581824 496108
rect 576597 495764 576965 495788
rect 579364 485722 581824 495788
rect 579364 483310 579388 485722
rect 581800 483310 581824 485722
rect 579364 448070 581824 483310
rect 579364 445658 579388 448070
rect 581800 445658 581824 448070
rect 579364 423070 581824 445658
rect 579175 422711 581824 423070
rect 578831 422687 581824 422711
rect 578831 422367 578855 422687
rect 579175 422367 581824 422687
rect 578831 422343 581824 422367
rect 579175 421791 581824 422343
rect 579364 417852 581824 421791
rect 579522 417032 581824 417852
rect 27813 416997 28663 417021
rect 27813 416195 27837 416997
rect 28639 416195 28663 416997
rect 27813 407398 28663 416195
rect 45037 407398 334930 415191
rect 578255 414750 578623 414774
rect 579364 414750 581824 417032
rect 578255 414430 578279 414750
rect 578599 414430 581824 414750
rect 578255 414406 578623 414430
rect 579364 409752 581824 414430
rect 5787 402491 6685 402515
rect 17306 402491 334930 407398
rect 5787 401641 5811 402491
rect 6661 401641 334930 402491
rect 5787 401617 6685 401641
rect 17306 398260 334930 401641
rect 45037 389569 334930 398260
rect 573026 407292 581824 409752
rect 573026 396574 575486 407292
rect 569970 396550 575486 396574
rect 569970 394138 569994 396550
rect 572406 394138 575486 396550
rect 569970 394114 575486 394138
rect 1698 336742 2538 336766
rect 1698 336414 1722 336742
rect 2050 336414 2538 336742
rect 1698 336390 2538 336414
rect 2162 303206 2538 336390
rect 259721 322855 287143 322879
rect 201547 307776 259745 322855
rect 2162 302830 6042 303206
rect 5666 242060 6042 302830
rect 201547 295481 204774 307776
rect 204750 293520 204774 295481
rect 219042 295481 259745 307776
rect 287119 295481 287143 322855
rect 219042 293520 219066 295481
rect 259721 295457 287143 295481
rect 204750 293496 219066 293520
rect 217578 287444 225148 287468
rect 109126 286274 112450 286298
rect 109126 285822 109150 286274
rect 109602 285822 112450 286274
rect 109126 285798 112450 285822
rect 110501 278490 110869 278514
rect 110501 278258 110525 278490
rect 110296 278170 110525 278258
rect 110845 278482 111236 278490
rect 111950 278482 112450 285798
rect 121208 285823 122866 285847
rect 126487 285823 131622 287187
rect 121208 284213 121232 285823
rect 122842 284213 131622 285823
rect 121208 284189 122866 284213
rect 110845 278170 112450 278482
rect 110296 277982 112450 278170
rect 110296 277860 111346 277982
rect 110267 277836 111346 277860
rect 110267 277516 110291 277836
rect 110611 277516 111346 277836
rect 110267 277492 111346 277516
rect 110272 277140 111346 277492
rect 110846 269208 111346 277140
rect 110846 269184 120326 269208
rect 110846 268732 119850 269184
rect 120302 268732 120326 269184
rect 110846 268708 120326 268732
rect 110846 268137 111346 268708
rect 110821 268113 111371 268137
rect 110821 267613 110845 268113
rect 111347 267613 111371 268113
rect 110821 267589 111371 267613
rect 126487 266868 131622 284213
rect 217578 279910 217602 287444
rect 225124 287438 225148 287444
rect 309308 287438 334930 389569
rect 225124 279916 334930 287438
rect 225124 279910 225148 279916
rect 217578 279886 225148 279910
rect 126487 266400 128674 266868
rect 129142 266400 131622 266868
rect 126487 263400 131622 266400
rect 126487 262932 128992 263400
rect 129460 262932 131622 263400
rect 88653 260951 89300 260959
rect 88653 260935 89640 260951
rect 88653 260653 88677 260935
rect 88959 260653 89640 260935
rect 88653 260629 89640 260653
rect 89013 260621 89640 260629
rect 87434 242066 87860 242090
rect 87434 242060 87458 242066
rect 5666 241684 87458 242060
rect 87434 241678 87458 241684
rect 87836 241678 87860 242066
rect 87434 241654 87860 241678
rect 89310 237192 89640 260621
rect 89182 236596 89936 237192
rect 89310 235033 89640 236596
rect 89280 235009 89670 235033
rect 89280 234679 89304 235009
rect 89646 234679 89670 235009
rect 89280 234655 89670 234679
rect 33238 231398 57778 233624
rect 33238 230762 35449 231398
rect 36083 230762 57778 231398
rect 33238 189802 57778 230762
rect 126487 221937 131622 262932
rect 309308 228238 334930 279916
rect 573026 288011 575486 394114
rect 573026 287691 573372 288011
rect 573692 287691 575486 288011
rect 573026 228238 575486 287691
rect 309308 227442 575486 228238
rect 306320 227156 575486 227442
rect 126487 216802 134198 221937
rect 129063 199264 134198 216802
rect 305406 221050 575486 227156
rect 305406 204923 581180 221050
rect 305406 204899 581205 204923
rect 305406 202616 558615 204899
rect 129036 199240 134224 199264
rect 129036 194100 129060 199240
rect 134200 194100 134224 199240
rect 129036 194076 134224 194100
rect 305406 189802 329946 202616
rect 33238 189778 329946 189802
rect 33238 184158 102584 189778
rect 108204 184158 329946 189778
rect 33238 157130 329946 184158
rect 558591 182335 558615 202616
rect 581181 182335 581205 204899
rect 558591 182311 581205 182335
<< comment >>
rect -100 704000 584100 704100
rect -100 0 0 704000
rect 584000 0 584100 704000
rect -100 -100 584100 0
use analogsub  analogsub_0 ~/caravel_user_project_analog/mag/./magicwrap/analogsub
timestamp 1672350823
transform 1 0 167268 0 1 254349
box -1480 -897 1606 3002
use analogsub  analogsub_1
timestamp 1672350823
transform 1 0 167284 0 1 247941
box -1480 -897 1606 3002
use analogsub  analogsub_2
timestamp 1672350823
transform 0 -1 15446 1 0 343536
box -1480 -897 1606 3002
use clkdiv  clkdiv_0 ~/caravel_user_project_analog/mag/./magicwrap/clkdiv
timestamp 1672477588
transform 0 -1 576260 1 0 410230
box 1566 -110 6170 3040
use filter  filter_0 ~/caravel_user_project_analog/mag/./magicwrap/filter
timestamp 1672466235
transform 1 0 155492 0 1 259112
box 17860 -47400 26372 -13499
use filter  filter_1
timestamp 1672466235
transform 1 0 165682 0 1 259002
box 17860 -47400 26372 -13499
use gilbert  gilbert_0 ~/caravel_user_project_analog/mag/./magicwrap/gilbert
timestamp 1672366060
transform 1 0 110361 0 1 273204
box -4331 -2998 105 2451
use gilbert  gilbert_1
timestamp 1672366060
transform 1 0 110415 0 1 282750
box -4331 -2998 105 2451
use opamp  opamp_0 ~/caravel_user_project_analog/mag/./magicwrap/opamp
timestamp 1672366615
transform 1 0 212190 0 1 287968
box -4400 -200 13580 6080
use opamp  opamp_1
timestamp 1672366615
transform 0 -1 10972 1 0 311798
box -4400 -200 13580 6080
use opamp  opamp_2
timestamp 1672366615
transform 0 -1 23232 1 0 414058
box -4400 -200 13580 6080
use phasecmp  phasecmp_0 ~/caravel_user_project_analog/mag/./magicwrap/phasecmp
timestamp 1672477588
transform 0 -1 576721 1 0 417218
box -1900 -2163 9838 -241
use quadgen  quadgen_0 ~/caravel_user_project_analog/mag/./magicwrap/quadgen
timestamp 1672477588
transform 1 0 104418 0 1 288480
box -428 -410 8928 644
use sky130_fd_pr__cap_mim_m3_1_2FRDLY  sky130_fd_pr__cap_mim_m3_1_2FRDLY_0
timestamp 1672468335
transform 1 0 580905 0 1 287351
box -1187 -1041 1187 1041
use sky130_fd_pr__cap_mim_m3_1_5B6GLN  sky130_fd_pr__cap_mim_m3_1_5B6GLN_0
timestamp 1672468335
transform 1 0 580759 0 1 297715
box -1687 -1541 1687 1541
use sky130_fd_pr__cap_mim_m3_1_P68BUM  sky130_fd_pr__cap_mim_m3_1_P68BUM_0
timestamp 1672468335
transform 1 0 41160 0 1 265138
box -3186 -3040 3186 3040
use sky130_fd_pr__cap_mim_m3_1_P68BUM  sky130_fd_pr__cap_mim_m3_1_P68BUM_1
timestamp 1672468335
transform 1 0 69098 0 1 282448
box -3186 -3040 3186 3040
use sky130_fd_pr__cap_mim_m3_1_P68BUM  sky130_fd_pr__cap_mim_m3_1_P68BUM_2
timestamp 1672468335
transform 1 0 20180 0 1 431712
box -3186 -3040 3186 3040
use sky130_fd_pr__cap_mim_m3_1_P68BUM  sky130_fd_pr__cap_mim_m3_1_P68BUM_3
timestamp 1672468335
transform 1 0 7362 0 1 333534
box -3186 -3040 3186 3040
use sky130_fd_pr__cap_mim_m3_1_P68BUM  sky130_fd_pr__cap_mim_m3_1_P68BUM_4
timestamp 1672468335
transform 1 0 8126 0 1 303630
box -3186 -3040 3186 3040
use sky130_fd_pr__cap_mim_m3_1_P68BUM  sky130_fd_pr__cap_mim_m3_1_P68BUM_5
timestamp 1672468335
transform 1 0 199232 0 1 286184
box -3186 -3040 3186 3040
use sky130_fd_pr__cap_mim_m3_1_PUMBUM  sky130_fd_pr__cap_mim_m3_1_PUMBUM_0
timestamp 1672468335
transform 1 0 20014 0 1 257158
box -13104 -12640 13104 12640
use sky130_fd_pr__cap_mim_m3_1_PUMBUM  sky130_fd_pr__cap_mim_m3_1_PUMBUM_1
timestamp 1672468335
transform 1 0 65168 0 1 253816
box -13104 -12640 13104 12640
use sky130_fd_pr__cap_mim_m3_1_PUMBUM  sky130_fd_pr__cap_mim_m3_1_PUMBUM_2
timestamp 1672468335
transform 1 0 52062 0 1 282430
box -13104 -12640 13104 12640
use sky130_fd_pr__cap_mim_m3_1_PUMBUM  sky130_fd_pr__cap_mim_m3_1_PUMBUM_3
timestamp 1672468335
transform 1 0 85858 0 1 282580
box -13104 -12640 13104 12640
use sky130_fd_pr__cap_mim_m3_1_PUMBUM  sky130_fd_pr__cap_mim_m3_1_PUMBUM_4
timestamp 1672468335
transform 1 0 106454 0 1 253568
box -13104 -12640 13104 12640
use sky130_fd_pr__cap_mim_m3_1_PUMBUM  sky130_fd_pr__cap_mim_m3_1_PUMBUM_5
timestamp 1672468335
transform 1 0 106122 0 1 225382
box -13104 -12640 13104 12640
use sky130_fd_pr__cap_mim_m3_1_PUMBUM  sky130_fd_pr__cap_mim_m3_1_PUMBUM_6
timestamp 1672468335
transform 1 0 146266 0 1 277490
box -13104 -12640 13104 12640
use sky130_fd_pr__cap_mim_m3_1_PUMBUM  sky130_fd_pr__cap_mim_m3_1_PUMBUM_7
timestamp 1672468335
transform 1 0 145904 0 1 248394
box -13104 -12640 13104 12640
use sky130_fd_pr__cap_mim_m3_1_PUMBUM  sky130_fd_pr__cap_mim_m3_1_PUMBUM_8
timestamp 1672468335
transform 1 0 145990 0 1 306504
box -13104 -12640 13104 12640
use sky130_fd_pr__cap_mim_m3_1_PUMBUM  sky130_fd_pr__cap_mim_m3_1_PUMBUM_9
timestamp 1672468335
transform 1 0 146094 0 1 336728
box -13104 -12640 13104 12640
use sky130_fd_pr__cap_mim_m3_1_PUMBUM  sky130_fd_pr__cap_mim_m3_1_PUMBUM_10
timestamp 1672468335
transform 1 0 23488 0 1 378116
box -13104 -12640 13104 12640
use sky130_fd_pr__cap_mim_m3_1_PUMBUM  sky130_fd_pr__cap_mim_m3_1_PUMBUM_11
timestamp 1672468335
transform 1 0 224650 0 1 259864
box -13104 -12640 13104 12640
use sky130_fd_pr__cap_mim_m3_1_PUMBUM  sky130_fd_pr__cap_mim_m3_1_PUMBUM_12
timestamp 1672468335
transform 1 0 224940 0 1 227676
box -13104 -12640 13104 12640
use sky130_fd_pr__cap_mim_m3_1_R8KP6D  sky130_fd_pr__cap_mim_m3_1_R8KP6D_0
timestamp 1672468335
transform 1 0 18904 0 1 322942
box -5454 -5282 5454 5282
use sky130_fd_pr__cap_mim_m3_1_REKGFF  sky130_fd_pr__cap_mim_m3_1_REKGFF_0
timestamp 1672474592
transform 1 0 40763 0 1 258631
box -2687 -2541 2687 2541
use sky130_fd_pr__cap_mim_m3_1_REKGFF  sky130_fd_pr__cap_mim_m3_1_REKGFF_1
timestamp 1672474592
transform 1 0 79093 0 1 231337
box -2687 -2541 2687 2541
use sky130_fd_pr__cap_mim_m3_1_REKGFF  sky130_fd_pr__cap_mim_m3_1_REKGFF_2
timestamp 1672474592
transform 1 0 116707 0 1 290789
box -2687 -2541 2687 2541
use sky130_fd_pr__cap_mim_m3_1_REKGFF  sky130_fd_pr__cap_mim_m3_1_REKGFF_3
timestamp 1672474592
transform 1 0 167417 0 1 242235
box -2687 -2541 2687 2541
use sky130_fd_pr__cap_mim_m3_1_REKGFF  sky130_fd_pr__cap_mim_m3_1_REKGFF_4
timestamp 1672474592
transform 1 0 173735 0 1 254693
box -2687 -2541 2687 2541
use sky130_fd_pr__cap_mim_m3_1_REKGFF  sky130_fd_pr__cap_mim_m3_1_REKGFF_5
timestamp 1672474592
transform -1 0 574255 0 -1 401993
box -2687 -2541 2687 2541
use sky130_fd_pr__cap_mim_m3_1_REKGFF  sky130_fd_pr__cap_mim_m3_1_REKGFF_6
timestamp 1672474592
transform 1 0 577453 0 1 452903
box -2687 -2541 2687 2541
use sky130_fd_pr__cap_mim_m3_1_REKGFF  sky130_fd_pr__cap_mim_m3_1_REKGFF_7
timestamp 1672474592
transform 1 0 576077 0 1 489969
box -2687 -2541 2687 2541
use sky130_fd_pr__nfet_01v8_JFBZSQ  sky130_fd_pr__nfet_01v8_JFBZSQ_0
timestamp 1672468335
transform 1 0 580498 0 1 292211
box -497 -2210 497 2210
use sky130_fd_pr__nfet_01v8_lvt_JDBWNB  sky130_fd_pr__nfet_01v8_lvt_JDBWNB_0
timestamp 1672468335
transform 1 0 36363 0 1 257287
box -246 -1210 246 1210
use sky130_fd_pr__nfet_01v8_lvt_U9BGXT  sky130_fd_pr__nfet_01v8_lvt_U9BGXT_0
timestamp 1672468335
transform 1 0 87169 0 1 251811
box -246 -510 246 510
use sky130_fd_pr__pfet_01v8_GXFJV8  sky130_fd_pr__pfet_01v8_GXFJV8_0
timestamp 1672468335
transform 1 0 579098 0 1 292219
box -497 -2219 497 2219
use sky130_fd_pr__pfet_01v8_lvt_3LXTS5  sky130_fd_pr__pfet_01v8_lvt_3LXTS5_0
timestamp 1672468335
transform 1 0 85807 0 1 255537
box -246 -519 246 519
use sky130_fd_pr__pfet_01v8_lvt_TDASS5  sky130_fd_pr__pfet_01v8_lvt_TDASS5_0
timestamp 1672468335
transform 1 0 35337 0 1 258029
box -246 -719 246 719
use sky130_fd_pr__pfet_01v8_lvt_TDASS5  sky130_fd_pr__pfet_01v8_lvt_TDASS5_1
timestamp 1672468335
transform 1 0 35337 0 1 259457
box -246 -719 246 719
use sky130_fd_pr__pfet_01v8_lvt_TRXTS5  sky130_fd_pr__pfet_01v8_lvt_TRXTS5_1
timestamp 1672468335
transform 1 0 36360 0 1 259380
box -246 -719 246 719
use sky130_fd_pr__pfet_01v8_lvt_XM7B29  sky130_fd_pr__pfet_01v8_lvt_XM7B29_0
timestamp 1672468335
transform 1 0 67956 0 1 277504
box -246 -1219 246 1219
use sky130_fd_pr__pfet_01v8_lvt_XRYC29  sky130_fd_pr__pfet_01v8_lvt_XRYC29_0
timestamp 1672468335
transform 1 0 67987 0 1 274627
box -246 -1219 246 1219
use sky130_fd_pr__res_xhigh_po_0p35_G3F5X4  sky130_fd_pr__res_xhigh_po_0p35_G3F5X4_0
timestamp 1672468335
transform 1 0 35097 0 1 267727
box -201 -3598 201 3598
use sky130_fd_pr__res_xhigh_po_0p35_G3F5X4  sky130_fd_pr__res_xhigh_po_0p35_G3F5X4_1
timestamp 1672468335
transform 1 0 87181 0 1 264045
box -201 -3598 201 3598
use sky130_fd_pr__res_xhigh_po_0p35_G3F5X4  sky130_fd_pr__res_xhigh_po_0p35_G3F5X4_2
timestamp 1672468335
transform 1 0 123195 0 1 240365
box -201 -3598 201 3598
use sky130_fd_pr__res_xhigh_po_0p35_G3F5X4  sky130_fd_pr__res_xhigh_po_0p35_G3F5X4_3
timestamp 1672468335
transform 1 0 124324 0 1 240316
box -201 -3598 201 3598
use sky130_fd_pr__res_xhigh_po_0p35_G3F5X4  sky130_fd_pr__res_xhigh_po_0p35_G3F5X4_4
timestamp 1672468335
transform 1 0 125344 0 1 240288
box -201 -3598 201 3598
use sky130_fd_pr__res_xhigh_po_0p35_G3F5X4  sky130_fd_pr__res_xhigh_po_0p35_G3F5X4_5
timestamp 1672468335
transform 1 0 126378 0 1 240282
box -201 -3598 201 3598
use sky130_fd_pr__res_xhigh_po_0p35_G3F5X4  sky130_fd_pr__res_xhigh_po_0p35_G3F5X4_6
timestamp 1672468335
transform 1 0 195175 0 1 217623
box -201 -3598 201 3598
use sky130_fd_pr__res_xhigh_po_0p35_G3F5X4  sky130_fd_pr__res_xhigh_po_0p35_G3F5X4_7
timestamp 1672468335
transform 1 0 197868 0 1 217642
box -201 -3598 201 3598
use sky130_fd_pr__res_xhigh_po_0p35_LU79P3  sky130_fd_pr__res_xhigh_po_0p35_LU79P3_0
timestamp 1672468335
transform 1 0 8321 0 1 326178
box -201 -1469 201 1469
use sky130_fd_pr__res_xhigh_po_0p35_LU79P3  sky130_fd_pr__res_xhigh_po_0p35_LU79P3_1
timestamp 1672468335
transform 0 1 9998 -1 0 327939
box -201 -1469 201 1469
use sky130_fd_pr__res_xhigh_po_0p35_R9FY7S  sky130_fd_pr__res_xhigh_po_0p35_R9FY7S_0
timestamp 1672468335
transform 1 0 87157 0 1 254414
box -201 -1649 201 1649
use sky130_fd_pr__res_xhigh_po_0p35_R9FY7S  sky130_fd_pr__res_xhigh_po_0p35_R9FY7S_1
timestamp 1672468335
transform 1 0 85779 0 1 252876
box -201 -1649 201 1649
use sky130_fd_pr__res_xhigh_po_0p35_ZSYV2F  sky130_fd_pr__res_xhigh_po_0p35_ZSYV2F_0
timestamp 1672468335
transform 1 0 9408 0 1 366695
box -201 -3599 201 3599
use sky130_fd_pr__res_xhigh_po_5p73_P7BAXV  sky130_fd_pr__res_xhigh_po_5p73_P7BAXV_0
timestamp 1672468335
transform 1 0 85095 0 1 234118
box -739 -1599 739 1599
use sky130_fd_pr__res_xhigh_po_5p73_P7BAXV  sky130_fd_pr__res_xhigh_po_5p73_P7BAXV_1
timestamp 1672468335
transform 1 0 85089 0 1 230460
box -739 -1599 739 1599
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1669390400
transform 1 0 579768 0 1 295218
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_1
timestamp 1669390400
transform 0 1 571314 -1 0 503246
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1669390400
transform 1 0 579584 0 1 295220
box -38 -48 130 592
use vco  vco_0 ~/caravel_user_project_analog/mag/./magicwrap/vco
timestamp 1672477588
transform 0 -1 574912 1 0 496541
box -2285 -199 4820 6220
<< labels >>
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1120 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s -800 381864 480 381976 0 FreeSans 1120 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s -800 338642 480 338754 0 FreeSans 1120 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -800 295420 480 295532 0 FreeSans 1120 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -800 252398 480 252510 0 FreeSans 1120 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s -800 124776 480 124888 0 FreeSans 1120 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s -800 81554 480 81666 0 FreeSans 1120 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s -800 38332 480 38444 0 FreeSans 1120 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -800 16910 480 17022 0 FreeSans 1120 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1120 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1120 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1120 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1120 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1120 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1120 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s -800 511530 480 511642 0 FreeSans 1120 0 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s -800 468308 480 468420 0 FreeSans 1120 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal3 s -800 425086 480 425198 0 FreeSans 1120 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1120 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s -800 380682 480 380794 0 FreeSans 1120 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s -800 337460 480 337572 0 FreeSans 1120 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s -800 294238 480 294350 0 FreeSans 1120 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -800 251216 480 251328 0 FreeSans 1120 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -800 123594 480 123706 0 FreeSans 1120 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -800 80372 480 80484 0 FreeSans 1120 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s -800 37150 480 37262 0 FreeSans 1120 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s -800 15728 480 15840 0 FreeSans 1120 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1120 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1120 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1120 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1120 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1120 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1120 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s -800 510348 480 510460 0 FreeSans 1120 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s -800 467126 480 467238 0 FreeSans 1120 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -800 423904 480 424016 0 FreeSans 1120 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1120 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1120 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 1920 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 1920 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 1920 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal4 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 1920 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 1920 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 1920 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 1920 180 0 0 io_clamp_high[0]
port 50 nsew signal bidirectional
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 1920 180 0 0 io_clamp_high[1]
port 51 nsew signal bidirectional
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 1920 180 0 0 io_clamp_high[2]
port 52 nsew signal bidirectional
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 1920 180 0 0 io_clamp_low[0]
port 53 nsew signal bidirectional
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 1920 180 0 0 io_clamp_low[1]
port 54 nsew signal bidirectional
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 1920 180 0 0 io_clamp_low[2]
port 55 nsew signal bidirectional
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1120 0 0 0 io_in[0]
port 56 nsew signal input
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1120 0 0 0 io_in[10]
port 57 nsew signal input
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1120 0 0 0 io_in[11]
port 58 nsew signal input
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1120 0 0 0 io_in[12]
port 59 nsew signal input
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1120 0 0 0 io_in[13]
port 60 nsew signal input
flabel metal3 s -800 507984 480 508096 0 FreeSans 1120 0 0 0 io_in[14]
port 61 nsew signal input
flabel metal3 s -800 464762 480 464874 0 FreeSans 1120 0 0 0 io_in[15]
port 62 nsew signal input
flabel metal3 s -800 421540 480 421652 0 FreeSans 1120 0 0 0 io_in[16]
port 63 nsew signal input
flabel metal3 s -800 378318 480 378430 0 FreeSans 1120 0 0 0 io_in[17]
port 64 nsew signal input
flabel metal3 s -800 335096 480 335208 0 FreeSans 1120 0 0 0 io_in[18]
port 65 nsew signal input
flabel metal3 s -800 291874 480 291986 0 FreeSans 1120 0 0 0 io_in[19]
port 66 nsew signal input
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1120 0 0 0 io_in[1]
port 67 nsew signal input
flabel metal3 s -800 248852 480 248964 0 FreeSans 1120 0 0 0 io_in[20]
port 68 nsew signal input
flabel metal3 s -800 121230 480 121342 0 FreeSans 1120 0 0 0 io_in[21]
port 69 nsew signal input
flabel metal3 s -800 78008 480 78120 0 FreeSans 1120 0 0 0 io_in[22]
port 70 nsew signal input
flabel metal3 s -800 34786 480 34898 0 FreeSans 1120 0 0 0 io_in[23]
port 71 nsew signal input
flabel metal3 s -800 13364 480 13476 0 FreeSans 1120 0 0 0 io_in[24]
port 72 nsew signal input
flabel metal3 s -800 8636 480 8748 0 FreeSans 1120 0 0 0 io_in[25]
port 73 nsew signal input
flabel metal3 s -800 3908 480 4020 0 FreeSans 1120 0 0 0 io_in[26]
port 74 nsew signal input
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1120 0 0 0 io_in[2]
port 75 nsew signal input
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1120 0 0 0 io_in[3]
port 76 nsew signal input
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1120 0 0 0 io_in[4]
port 77 nsew signal input
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1120 0 0 0 io_in[5]
port 78 nsew signal input
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1120 0 0 0 io_in[6]
port 79 nsew signal input
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1120 0 0 0 io_in[7]
port 80 nsew signal input
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1120 0 0 0 io_in[8]
port 81 nsew signal input
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1120 0 0 0 io_in[9]
port 82 nsew signal input
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1120 0 0 0 io_in_3v3[0]
port 83 nsew signal input
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1120 0 0 0 io_in_3v3[10]
port 84 nsew signal input
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1120 0 0 0 io_in_3v3[11]
port 85 nsew signal input
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1120 0 0 0 io_in_3v3[12]
port 86 nsew signal input
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1120 0 0 0 io_in_3v3[13]
port 87 nsew signal input
flabel metal3 s -800 509166 480 509278 0 FreeSans 1120 0 0 0 io_in_3v3[14]
port 88 nsew signal input
flabel metal3 s -800 465944 480 466056 0 FreeSans 1120 0 0 0 io_in_3v3[15]
port 89 nsew signal input
flabel metal3 s -800 422722 480 422834 0 FreeSans 1120 0 0 0 io_in_3v3[16]
port 90 nsew signal input
flabel metal3 s -800 379500 480 379612 0 FreeSans 1120 0 0 0 io_in_3v3[17]
port 91 nsew signal input
flabel metal3 s -800 336278 480 336390 0 FreeSans 1120 0 0 0 io_in_3v3[18]
port 92 nsew signal input
flabel metal3 s -800 293056 480 293168 0 FreeSans 1120 0 0 0 io_in_3v3[19]
port 93 nsew signal input
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1120 0 0 0 io_in_3v3[1]
port 94 nsew signal input
flabel metal3 s -800 250034 480 250146 0 FreeSans 1120 0 0 0 io_in_3v3[20]
port 95 nsew signal input
flabel metal3 s -800 122412 480 122524 0 FreeSans 1120 0 0 0 io_in_3v3[21]
port 96 nsew signal input
flabel metal3 s -800 79190 480 79302 0 FreeSans 1120 0 0 0 io_in_3v3[22]
port 97 nsew signal input
flabel metal3 s -800 35968 480 36080 0 FreeSans 1120 0 0 0 io_in_3v3[23]
port 98 nsew signal input
flabel metal3 s -800 14546 480 14658 0 FreeSans 1120 0 0 0 io_in_3v3[24]
port 99 nsew signal input
flabel metal3 s -800 9818 480 9930 0 FreeSans 1120 0 0 0 io_in_3v3[25]
port 100 nsew signal input
flabel metal3 s -800 5090 480 5202 0 FreeSans 1120 0 0 0 io_in_3v3[26]
port 101 nsew signal input
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1120 0 0 0 io_in_3v3[2]
port 102 nsew signal input
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1120 0 0 0 io_in_3v3[3]
port 103 nsew signal input
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1120 0 0 0 io_in_3v3[4]
port 104 nsew signal input
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1120 0 0 0 io_in_3v3[5]
port 105 nsew signal input
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1120 0 0 0 io_in_3v3[6]
port 106 nsew signal input
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1120 0 0 0 io_in_3v3[7]
port 107 nsew signal input
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1120 0 0 0 io_in_3v3[8]
port 108 nsew signal input
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1120 0 0 0 io_in_3v3[9]
port 109 nsew signal input
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1120 0 0 0 io_oeb[0]
port 110 nsew signal tristate
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1120 0 0 0 io_oeb[10]
port 111 nsew signal tristate
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1120 0 0 0 io_oeb[11]
port 112 nsew signal tristate
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1120 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1120 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s -800 505620 480 505732 0 FreeSans 1120 0 0 0 io_oeb[14]
port 115 nsew signal tristate
flabel metal3 s -800 462398 480 462510 0 FreeSans 1120 0 0 0 io_oeb[15]
port 116 nsew signal tristate
flabel metal3 s -800 419176 480 419288 0 FreeSans 1120 0 0 0 io_oeb[16]
port 117 nsew signal tristate
flabel metal3 s -800 375954 480 376066 0 FreeSans 1120 0 0 0 io_oeb[17]
port 118 nsew signal tristate
flabel metal3 s -800 332732 480 332844 0 FreeSans 1120 0 0 0 io_oeb[18]
port 119 nsew signal tristate
flabel metal3 s -800 289510 480 289622 0 FreeSans 1120 0 0 0 io_oeb[19]
port 120 nsew signal tristate
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1120 0 0 0 io_oeb[1]
port 121 nsew signal tristate
flabel metal3 s -800 246488 480 246600 0 FreeSans 1120 0 0 0 io_oeb[20]
port 122 nsew signal tristate
flabel metal3 s -800 118866 480 118978 0 FreeSans 1120 0 0 0 io_oeb[21]
port 123 nsew signal tristate
flabel metal3 s -800 75644 480 75756 0 FreeSans 1120 0 0 0 io_oeb[22]
port 124 nsew signal tristate
flabel metal3 s -800 32422 480 32534 0 FreeSans 1120 0 0 0 io_oeb[23]
port 125 nsew signal tristate
flabel metal3 s -800 11000 480 11112 0 FreeSans 1120 0 0 0 io_oeb[24]
port 126 nsew signal tristate
flabel metal3 s -800 6272 480 6384 0 FreeSans 1120 0 0 0 io_oeb[25]
port 127 nsew signal tristate
flabel metal3 s -800 1544 480 1656 0 FreeSans 1120 0 0 0 io_oeb[26]
port 128 nsew signal tristate
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1120 0 0 0 io_oeb[2]
port 129 nsew signal tristate
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1120 0 0 0 io_oeb[3]
port 130 nsew signal tristate
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1120 0 0 0 io_oeb[4]
port 131 nsew signal tristate
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1120 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1120 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1120 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1120 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1120 0 0 0 io_oeb[9]
port 136 nsew signal tristate
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1120 0 0 0 io_out[0]
port 137 nsew signal tristate
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1120 0 0 0 io_out[10]
port 138 nsew signal tristate
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1120 0 0 0 io_out[11]
port 139 nsew signal tristate
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1120 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1120 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s -800 506802 480 506914 0 FreeSans 1120 0 0 0 io_out[14]
port 142 nsew signal tristate
flabel metal3 s -800 463580 480 463692 0 FreeSans 1120 0 0 0 io_out[15]
port 143 nsew signal tristate
flabel metal3 s -800 420358 480 420470 0 FreeSans 1120 0 0 0 io_out[16]
port 144 nsew signal tristate
flabel metal3 s -800 377136 480 377248 0 FreeSans 1120 0 0 0 io_out[17]
port 145 nsew signal tristate
flabel metal3 s -800 333914 480 334026 0 FreeSans 1120 0 0 0 io_out[18]
port 146 nsew signal tristate
flabel metal3 s -800 290692 480 290804 0 FreeSans 1120 0 0 0 io_out[19]
port 147 nsew signal tristate
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1120 0 0 0 io_out[1]
port 148 nsew signal tristate
flabel metal3 s -800 247670 480 247782 0 FreeSans 1120 0 0 0 io_out[20]
port 149 nsew signal tristate
flabel metal3 s -800 120048 480 120160 0 FreeSans 1120 0 0 0 io_out[21]
port 150 nsew signal tristate
flabel metal3 s -800 76826 480 76938 0 FreeSans 1120 0 0 0 io_out[22]
port 151 nsew signal tristate
flabel metal3 s -800 33604 480 33716 0 FreeSans 1120 0 0 0 io_out[23]
port 152 nsew signal tristate
flabel metal3 s -800 12182 480 12294 0 FreeSans 1120 0 0 0 io_out[24]
port 153 nsew signal tristate
flabel metal3 s -800 7454 480 7566 0 FreeSans 1120 0 0 0 io_out[25]
port 154 nsew signal tristate
flabel metal3 s -800 2726 480 2838 0 FreeSans 1120 0 0 0 io_out[26]
port 155 nsew signal tristate
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1120 0 0 0 io_out[2]
port 156 nsew signal tristate
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1120 0 0 0 io_out[3]
port 157 nsew signal tristate
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1120 0 0 0 io_out[4]
port 158 nsew signal tristate
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1120 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1120 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1120 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1120 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1120 0 0 0 io_out[9]
port 163 nsew signal tristate
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1120 90 0 0 la_data_in[0]
port 164 nsew signal input
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1120 90 0 0 la_data_in[100]
port 165 nsew signal input
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1120 90 0 0 la_data_in[101]
port 166 nsew signal input
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1120 90 0 0 la_data_in[102]
port 167 nsew signal input
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1120 90 0 0 la_data_in[103]
port 168 nsew signal input
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1120 90 0 0 la_data_in[104]
port 169 nsew signal input
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1120 90 0 0 la_data_in[105]
port 170 nsew signal input
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1120 90 0 0 la_data_in[106]
port 171 nsew signal input
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1120 90 0 0 la_data_in[107]
port 172 nsew signal input
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1120 90 0 0 la_data_in[108]
port 173 nsew signal input
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1120 90 0 0 la_data_in[109]
port 174 nsew signal input
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1120 90 0 0 la_data_in[10]
port 175 nsew signal input
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1120 90 0 0 la_data_in[110]
port 176 nsew signal input
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1120 90 0 0 la_data_in[111]
port 177 nsew signal input
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1120 90 0 0 la_data_in[112]
port 178 nsew signal input
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1120 90 0 0 la_data_in[113]
port 179 nsew signal input
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1120 90 0 0 la_data_in[114]
port 180 nsew signal input
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1120 90 0 0 la_data_in[115]
port 181 nsew signal input
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1120 90 0 0 la_data_in[116]
port 182 nsew signal input
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1120 90 0 0 la_data_in[117]
port 183 nsew signal input
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1120 90 0 0 la_data_in[118]
port 184 nsew signal input
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1120 90 0 0 la_data_in[119]
port 185 nsew signal input
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1120 90 0 0 la_data_in[11]
port 186 nsew signal input
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1120 90 0 0 la_data_in[120]
port 187 nsew signal input
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1120 90 0 0 la_data_in[121]
port 188 nsew signal input
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1120 90 0 0 la_data_in[122]
port 189 nsew signal input
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1120 90 0 0 la_data_in[123]
port 190 nsew signal input
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1120 90 0 0 la_data_in[124]
port 191 nsew signal input
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1120 90 0 0 la_data_in[125]
port 192 nsew signal input
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1120 90 0 0 la_data_in[126]
port 193 nsew signal input
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1120 90 0 0 la_data_in[127]
port 194 nsew signal input
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1120 90 0 0 la_data_in[12]
port 195 nsew signal input
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1120 90 0 0 la_data_in[13]
port 196 nsew signal input
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1120 90 0 0 la_data_in[14]
port 197 nsew signal input
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1120 90 0 0 la_data_in[15]
port 198 nsew signal input
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1120 90 0 0 la_data_in[16]
port 199 nsew signal input
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1120 90 0 0 la_data_in[17]
port 200 nsew signal input
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1120 90 0 0 la_data_in[18]
port 201 nsew signal input
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1120 90 0 0 la_data_in[19]
port 202 nsew signal input
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1120 90 0 0 la_data_in[1]
port 203 nsew signal input
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1120 90 0 0 la_data_in[20]
port 204 nsew signal input
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1120 90 0 0 la_data_in[21]
port 205 nsew signal input
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1120 90 0 0 la_data_in[22]
port 206 nsew signal input
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1120 90 0 0 la_data_in[23]
port 207 nsew signal input
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1120 90 0 0 la_data_in[24]
port 208 nsew signal input
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1120 90 0 0 la_data_in[25]
port 209 nsew signal input
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1120 90 0 0 la_data_in[26]
port 210 nsew signal input
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1120 90 0 0 la_data_in[27]
port 211 nsew signal input
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1120 90 0 0 la_data_in[28]
port 212 nsew signal input
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1120 90 0 0 la_data_in[29]
port 213 nsew signal input
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1120 90 0 0 la_data_in[2]
port 214 nsew signal input
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1120 90 0 0 la_data_in[30]
port 215 nsew signal input
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1120 90 0 0 la_data_in[31]
port 216 nsew signal input
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1120 90 0 0 la_data_in[32]
port 217 nsew signal input
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1120 90 0 0 la_data_in[33]
port 218 nsew signal input
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1120 90 0 0 la_data_in[34]
port 219 nsew signal input
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1120 90 0 0 la_data_in[35]
port 220 nsew signal input
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1120 90 0 0 la_data_in[36]
port 221 nsew signal input
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1120 90 0 0 la_data_in[37]
port 222 nsew signal input
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1120 90 0 0 la_data_in[38]
port 223 nsew signal input
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1120 90 0 0 la_data_in[39]
port 224 nsew signal input
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1120 90 0 0 la_data_in[3]
port 225 nsew signal input
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1120 90 0 0 la_data_in[40]
port 226 nsew signal input
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1120 90 0 0 la_data_in[41]
port 227 nsew signal input
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1120 90 0 0 la_data_in[42]
port 228 nsew signal input
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1120 90 0 0 la_data_in[43]
port 229 nsew signal input
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1120 90 0 0 la_data_in[44]
port 230 nsew signal input
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1120 90 0 0 la_data_in[45]
port 231 nsew signal input
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1120 90 0 0 la_data_in[46]
port 232 nsew signal input
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1120 90 0 0 la_data_in[47]
port 233 nsew signal input
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1120 90 0 0 la_data_in[48]
port 234 nsew signal input
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1120 90 0 0 la_data_in[49]
port 235 nsew signal input
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1120 90 0 0 la_data_in[4]
port 236 nsew signal input
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1120 90 0 0 la_data_in[50]
port 237 nsew signal input
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1120 90 0 0 la_data_in[51]
port 238 nsew signal input
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1120 90 0 0 la_data_in[52]
port 239 nsew signal input
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1120 90 0 0 la_data_in[53]
port 240 nsew signal input
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1120 90 0 0 la_data_in[54]
port 241 nsew signal input
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1120 90 0 0 la_data_in[55]
port 242 nsew signal input
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1120 90 0 0 la_data_in[56]
port 243 nsew signal input
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1120 90 0 0 la_data_in[57]
port 244 nsew signal input
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1120 90 0 0 la_data_in[58]
port 245 nsew signal input
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1120 90 0 0 la_data_in[59]
port 246 nsew signal input
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1120 90 0 0 la_data_in[5]
port 247 nsew signal input
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1120 90 0 0 la_data_in[60]
port 248 nsew signal input
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1120 90 0 0 la_data_in[61]
port 249 nsew signal input
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1120 90 0 0 la_data_in[62]
port 250 nsew signal input
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1120 90 0 0 la_data_in[63]
port 251 nsew signal input
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1120 90 0 0 la_data_in[64]
port 252 nsew signal input
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1120 90 0 0 la_data_in[65]
port 253 nsew signal input
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1120 90 0 0 la_data_in[66]
port 254 nsew signal input
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1120 90 0 0 la_data_in[67]
port 255 nsew signal input
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1120 90 0 0 la_data_in[68]
port 256 nsew signal input
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1120 90 0 0 la_data_in[69]
port 257 nsew signal input
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1120 90 0 0 la_data_in[6]
port 258 nsew signal input
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1120 90 0 0 la_data_in[70]
port 259 nsew signal input
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1120 90 0 0 la_data_in[71]
port 260 nsew signal input
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1120 90 0 0 la_data_in[72]
port 261 nsew signal input
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1120 90 0 0 la_data_in[73]
port 262 nsew signal input
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1120 90 0 0 la_data_in[74]
port 263 nsew signal input
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1120 90 0 0 la_data_in[75]
port 264 nsew signal input
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1120 90 0 0 la_data_in[76]
port 265 nsew signal input
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1120 90 0 0 la_data_in[77]
port 266 nsew signal input
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1120 90 0 0 la_data_in[78]
port 267 nsew signal input
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1120 90 0 0 la_data_in[79]
port 268 nsew signal input
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1120 90 0 0 la_data_in[7]
port 269 nsew signal input
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1120 90 0 0 la_data_in[80]
port 270 nsew signal input
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1120 90 0 0 la_data_in[81]
port 271 nsew signal input
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1120 90 0 0 la_data_in[82]
port 272 nsew signal input
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1120 90 0 0 la_data_in[83]
port 273 nsew signal input
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1120 90 0 0 la_data_in[84]
port 274 nsew signal input
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1120 90 0 0 la_data_in[85]
port 275 nsew signal input
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1120 90 0 0 la_data_in[86]
port 276 nsew signal input
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1120 90 0 0 la_data_in[87]
port 277 nsew signal input
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1120 90 0 0 la_data_in[88]
port 278 nsew signal input
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1120 90 0 0 la_data_in[89]
port 279 nsew signal input
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1120 90 0 0 la_data_in[8]
port 280 nsew signal input
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1120 90 0 0 la_data_in[90]
port 281 nsew signal input
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1120 90 0 0 la_data_in[91]
port 282 nsew signal input
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1120 90 0 0 la_data_in[92]
port 283 nsew signal input
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1120 90 0 0 la_data_in[93]
port 284 nsew signal input
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1120 90 0 0 la_data_in[94]
port 285 nsew signal input
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1120 90 0 0 la_data_in[95]
port 286 nsew signal input
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1120 90 0 0 la_data_in[96]
port 287 nsew signal input
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1120 90 0 0 la_data_in[97]
port 288 nsew signal input
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1120 90 0 0 la_data_in[98]
port 289 nsew signal input
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1120 90 0 0 la_data_in[99]
port 290 nsew signal input
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1120 90 0 0 la_data_in[9]
port 291 nsew signal input
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1120 90 0 0 la_data_out[0]
port 292 nsew signal tristate
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1120 90 0 0 la_data_out[100]
port 293 nsew signal tristate
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1120 90 0 0 la_data_out[101]
port 294 nsew signal tristate
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1120 90 0 0 la_data_out[102]
port 295 nsew signal tristate
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1120 90 0 0 la_data_out[103]
port 296 nsew signal tristate
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1120 90 0 0 la_data_out[104]
port 297 nsew signal tristate
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1120 90 0 0 la_data_out[105]
port 298 nsew signal tristate
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1120 90 0 0 la_data_out[106]
port 299 nsew signal tristate
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1120 90 0 0 la_data_out[107]
port 300 nsew signal tristate
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1120 90 0 0 la_data_out[108]
port 301 nsew signal tristate
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1120 90 0 0 la_data_out[109]
port 302 nsew signal tristate
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1120 90 0 0 la_data_out[10]
port 303 nsew signal tristate
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1120 90 0 0 la_data_out[110]
port 304 nsew signal tristate
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1120 90 0 0 la_data_out[111]
port 305 nsew signal tristate
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1120 90 0 0 la_data_out[112]
port 306 nsew signal tristate
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1120 90 0 0 la_data_out[113]
port 307 nsew signal tristate
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1120 90 0 0 la_data_out[114]
port 308 nsew signal tristate
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1120 90 0 0 la_data_out[115]
port 309 nsew signal tristate
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1120 90 0 0 la_data_out[116]
port 310 nsew signal tristate
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1120 90 0 0 la_data_out[117]
port 311 nsew signal tristate
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1120 90 0 0 la_data_out[118]
port 312 nsew signal tristate
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1120 90 0 0 la_data_out[119]
port 313 nsew signal tristate
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1120 90 0 0 la_data_out[11]
port 314 nsew signal tristate
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1120 90 0 0 la_data_out[120]
port 315 nsew signal tristate
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1120 90 0 0 la_data_out[121]
port 316 nsew signal tristate
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1120 90 0 0 la_data_out[122]
port 317 nsew signal tristate
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1120 90 0 0 la_data_out[123]
port 318 nsew signal tristate
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1120 90 0 0 la_data_out[124]
port 319 nsew signal tristate
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1120 90 0 0 la_data_out[125]
port 320 nsew signal tristate
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1120 90 0 0 la_data_out[126]
port 321 nsew signal tristate
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1120 90 0 0 la_data_out[127]
port 322 nsew signal tristate
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1120 90 0 0 la_data_out[12]
port 323 nsew signal tristate
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1120 90 0 0 la_data_out[13]
port 324 nsew signal tristate
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1120 90 0 0 la_data_out[14]
port 325 nsew signal tristate
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1120 90 0 0 la_data_out[15]
port 326 nsew signal tristate
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1120 90 0 0 la_data_out[16]
port 327 nsew signal tristate
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1120 90 0 0 la_data_out[17]
port 328 nsew signal tristate
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1120 90 0 0 la_data_out[18]
port 329 nsew signal tristate
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1120 90 0 0 la_data_out[19]
port 330 nsew signal tristate
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1120 90 0 0 la_data_out[1]
port 331 nsew signal tristate
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1120 90 0 0 la_data_out[20]
port 332 nsew signal tristate
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1120 90 0 0 la_data_out[21]
port 333 nsew signal tristate
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1120 90 0 0 la_data_out[22]
port 334 nsew signal tristate
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1120 90 0 0 la_data_out[23]
port 335 nsew signal tristate
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1120 90 0 0 la_data_out[24]
port 336 nsew signal tristate
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1120 90 0 0 la_data_out[25]
port 337 nsew signal tristate
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1120 90 0 0 la_data_out[26]
port 338 nsew signal tristate
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1120 90 0 0 la_data_out[27]
port 339 nsew signal tristate
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1120 90 0 0 la_data_out[28]
port 340 nsew signal tristate
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1120 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1120 90 0 0 la_data_out[2]
port 342 nsew signal tristate
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1120 90 0 0 la_data_out[30]
port 343 nsew signal tristate
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1120 90 0 0 la_data_out[31]
port 344 nsew signal tristate
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1120 90 0 0 la_data_out[32]
port 345 nsew signal tristate
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1120 90 0 0 la_data_out[33]
port 346 nsew signal tristate
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1120 90 0 0 la_data_out[34]
port 347 nsew signal tristate
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1120 90 0 0 la_data_out[35]
port 348 nsew signal tristate
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1120 90 0 0 la_data_out[36]
port 349 nsew signal tristate
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1120 90 0 0 la_data_out[37]
port 350 nsew signal tristate
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1120 90 0 0 la_data_out[38]
port 351 nsew signal tristate
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1120 90 0 0 la_data_out[39]
port 352 nsew signal tristate
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1120 90 0 0 la_data_out[3]
port 353 nsew signal tristate
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1120 90 0 0 la_data_out[40]
port 354 nsew signal tristate
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1120 90 0 0 la_data_out[41]
port 355 nsew signal tristate
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1120 90 0 0 la_data_out[42]
port 356 nsew signal tristate
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1120 90 0 0 la_data_out[43]
port 357 nsew signal tristate
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1120 90 0 0 la_data_out[44]
port 358 nsew signal tristate
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1120 90 0 0 la_data_out[45]
port 359 nsew signal tristate
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1120 90 0 0 la_data_out[46]
port 360 nsew signal tristate
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1120 90 0 0 la_data_out[47]
port 361 nsew signal tristate
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1120 90 0 0 la_data_out[48]
port 362 nsew signal tristate
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1120 90 0 0 la_data_out[49]
port 363 nsew signal tristate
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1120 90 0 0 la_data_out[4]
port 364 nsew signal tristate
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1120 90 0 0 la_data_out[50]
port 365 nsew signal tristate
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1120 90 0 0 la_data_out[51]
port 366 nsew signal tristate
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1120 90 0 0 la_data_out[52]
port 367 nsew signal tristate
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1120 90 0 0 la_data_out[53]
port 368 nsew signal tristate
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1120 90 0 0 la_data_out[54]
port 369 nsew signal tristate
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1120 90 0 0 la_data_out[55]
port 370 nsew signal tristate
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1120 90 0 0 la_data_out[56]
port 371 nsew signal tristate
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1120 90 0 0 la_data_out[57]
port 372 nsew signal tristate
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1120 90 0 0 la_data_out[58]
port 373 nsew signal tristate
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1120 90 0 0 la_data_out[59]
port 374 nsew signal tristate
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1120 90 0 0 la_data_out[5]
port 375 nsew signal tristate
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1120 90 0 0 la_data_out[60]
port 376 nsew signal tristate
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1120 90 0 0 la_data_out[61]
port 377 nsew signal tristate
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1120 90 0 0 la_data_out[62]
port 378 nsew signal tristate
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1120 90 0 0 la_data_out[63]
port 379 nsew signal tristate
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1120 90 0 0 la_data_out[64]
port 380 nsew signal tristate
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1120 90 0 0 la_data_out[65]
port 381 nsew signal tristate
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1120 90 0 0 la_data_out[66]
port 382 nsew signal tristate
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1120 90 0 0 la_data_out[67]
port 383 nsew signal tristate
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1120 90 0 0 la_data_out[68]
port 384 nsew signal tristate
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1120 90 0 0 la_data_out[69]
port 385 nsew signal tristate
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1120 90 0 0 la_data_out[6]
port 386 nsew signal tristate
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1120 90 0 0 la_data_out[70]
port 387 nsew signal tristate
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1120 90 0 0 la_data_out[71]
port 388 nsew signal tristate
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1120 90 0 0 la_data_out[72]
port 389 nsew signal tristate
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1120 90 0 0 la_data_out[73]
port 390 nsew signal tristate
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1120 90 0 0 la_data_out[74]
port 391 nsew signal tristate
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1120 90 0 0 la_data_out[75]
port 392 nsew signal tristate
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1120 90 0 0 la_data_out[76]
port 393 nsew signal tristate
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1120 90 0 0 la_data_out[77]
port 394 nsew signal tristate
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1120 90 0 0 la_data_out[78]
port 395 nsew signal tristate
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1120 90 0 0 la_data_out[79]
port 396 nsew signal tristate
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1120 90 0 0 la_data_out[7]
port 397 nsew signal tristate
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1120 90 0 0 la_data_out[80]
port 398 nsew signal tristate
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1120 90 0 0 la_data_out[81]
port 399 nsew signal tristate
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1120 90 0 0 la_data_out[82]
port 400 nsew signal tristate
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1120 90 0 0 la_data_out[83]
port 401 nsew signal tristate
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1120 90 0 0 la_data_out[84]
port 402 nsew signal tristate
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1120 90 0 0 la_data_out[85]
port 403 nsew signal tristate
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1120 90 0 0 la_data_out[86]
port 404 nsew signal tristate
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1120 90 0 0 la_data_out[87]
port 405 nsew signal tristate
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1120 90 0 0 la_data_out[88]
port 406 nsew signal tristate
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1120 90 0 0 la_data_out[89]
port 407 nsew signal tristate
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1120 90 0 0 la_data_out[8]
port 408 nsew signal tristate
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1120 90 0 0 la_data_out[90]
port 409 nsew signal tristate
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1120 90 0 0 la_data_out[91]
port 410 nsew signal tristate
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1120 90 0 0 la_data_out[92]
port 411 nsew signal tristate
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1120 90 0 0 la_data_out[93]
port 412 nsew signal tristate
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1120 90 0 0 la_data_out[94]
port 413 nsew signal tristate
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1120 90 0 0 la_data_out[95]
port 414 nsew signal tristate
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1120 90 0 0 la_data_out[96]
port 415 nsew signal tristate
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1120 90 0 0 la_data_out[97]
port 416 nsew signal tristate
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1120 90 0 0 la_data_out[98]
port 417 nsew signal tristate
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1120 90 0 0 la_data_out[99]
port 418 nsew signal tristate
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1120 90 0 0 la_data_out[9]
port 419 nsew signal tristate
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1120 90 0 0 la_oenb[0]
port 420 nsew signal input
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1120 90 0 0 la_oenb[100]
port 421 nsew signal input
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1120 90 0 0 la_oenb[101]
port 422 nsew signal input
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1120 90 0 0 la_oenb[102]
port 423 nsew signal input
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1120 90 0 0 la_oenb[103]
port 424 nsew signal input
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1120 90 0 0 la_oenb[104]
port 425 nsew signal input
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1120 90 0 0 la_oenb[105]
port 426 nsew signal input
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1120 90 0 0 la_oenb[106]
port 427 nsew signal input
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1120 90 0 0 la_oenb[107]
port 428 nsew signal input
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1120 90 0 0 la_oenb[108]
port 429 nsew signal input
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1120 90 0 0 la_oenb[109]
port 430 nsew signal input
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1120 90 0 0 la_oenb[10]
port 431 nsew signal input
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1120 90 0 0 la_oenb[110]
port 432 nsew signal input
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1120 90 0 0 la_oenb[111]
port 433 nsew signal input
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1120 90 0 0 la_oenb[112]
port 434 nsew signal input
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1120 90 0 0 la_oenb[113]
port 435 nsew signal input
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1120 90 0 0 la_oenb[114]
port 436 nsew signal input
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1120 90 0 0 la_oenb[115]
port 437 nsew signal input
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1120 90 0 0 la_oenb[116]
port 438 nsew signal input
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1120 90 0 0 la_oenb[117]
port 439 nsew signal input
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1120 90 0 0 la_oenb[118]
port 440 nsew signal input
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1120 90 0 0 la_oenb[119]
port 441 nsew signal input
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1120 90 0 0 la_oenb[11]
port 442 nsew signal input
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1120 90 0 0 la_oenb[120]
port 443 nsew signal input
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1120 90 0 0 la_oenb[121]
port 444 nsew signal input
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1120 90 0 0 la_oenb[122]
port 445 nsew signal input
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1120 90 0 0 la_oenb[123]
port 446 nsew signal input
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1120 90 0 0 la_oenb[124]
port 447 nsew signal input
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1120 90 0 0 la_oenb[125]
port 448 nsew signal input
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1120 90 0 0 la_oenb[126]
port 449 nsew signal input
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1120 90 0 0 la_oenb[127]
port 450 nsew signal input
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1120 90 0 0 la_oenb[12]
port 451 nsew signal input
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1120 90 0 0 la_oenb[13]
port 452 nsew signal input
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1120 90 0 0 la_oenb[14]
port 453 nsew signal input
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1120 90 0 0 la_oenb[15]
port 454 nsew signal input
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1120 90 0 0 la_oenb[16]
port 455 nsew signal input
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1120 90 0 0 la_oenb[17]
port 456 nsew signal input
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1120 90 0 0 la_oenb[18]
port 457 nsew signal input
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1120 90 0 0 la_oenb[19]
port 458 nsew signal input
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1120 90 0 0 la_oenb[1]
port 459 nsew signal input
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1120 90 0 0 la_oenb[20]
port 460 nsew signal input
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1120 90 0 0 la_oenb[21]
port 461 nsew signal input
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1120 90 0 0 la_oenb[22]
port 462 nsew signal input
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1120 90 0 0 la_oenb[23]
port 463 nsew signal input
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1120 90 0 0 la_oenb[24]
port 464 nsew signal input
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1120 90 0 0 la_oenb[25]
port 465 nsew signal input
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1120 90 0 0 la_oenb[26]
port 466 nsew signal input
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1120 90 0 0 la_oenb[27]
port 467 nsew signal input
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1120 90 0 0 la_oenb[28]
port 468 nsew signal input
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1120 90 0 0 la_oenb[29]
port 469 nsew signal input
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1120 90 0 0 la_oenb[2]
port 470 nsew signal input
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1120 90 0 0 la_oenb[30]
port 471 nsew signal input
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1120 90 0 0 la_oenb[31]
port 472 nsew signal input
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1120 90 0 0 la_oenb[32]
port 473 nsew signal input
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1120 90 0 0 la_oenb[33]
port 474 nsew signal input
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1120 90 0 0 la_oenb[34]
port 475 nsew signal input
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1120 90 0 0 la_oenb[35]
port 476 nsew signal input
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1120 90 0 0 la_oenb[36]
port 477 nsew signal input
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1120 90 0 0 la_oenb[37]
port 478 nsew signal input
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1120 90 0 0 la_oenb[38]
port 479 nsew signal input
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1120 90 0 0 la_oenb[39]
port 480 nsew signal input
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1120 90 0 0 la_oenb[3]
port 481 nsew signal input
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1120 90 0 0 la_oenb[40]
port 482 nsew signal input
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1120 90 0 0 la_oenb[41]
port 483 nsew signal input
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1120 90 0 0 la_oenb[42]
port 484 nsew signal input
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1120 90 0 0 la_oenb[43]
port 485 nsew signal input
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1120 90 0 0 la_oenb[44]
port 486 nsew signal input
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1120 90 0 0 la_oenb[45]
port 487 nsew signal input
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1120 90 0 0 la_oenb[46]
port 488 nsew signal input
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1120 90 0 0 la_oenb[47]
port 489 nsew signal input
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1120 90 0 0 la_oenb[48]
port 490 nsew signal input
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1120 90 0 0 la_oenb[49]
port 491 nsew signal input
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1120 90 0 0 la_oenb[4]
port 492 nsew signal input
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1120 90 0 0 la_oenb[50]
port 493 nsew signal input
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1120 90 0 0 la_oenb[51]
port 494 nsew signal input
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1120 90 0 0 la_oenb[52]
port 495 nsew signal input
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1120 90 0 0 la_oenb[53]
port 496 nsew signal input
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1120 90 0 0 la_oenb[54]
port 497 nsew signal input
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1120 90 0 0 la_oenb[55]
port 498 nsew signal input
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1120 90 0 0 la_oenb[56]
port 499 nsew signal input
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1120 90 0 0 la_oenb[57]
port 500 nsew signal input
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1120 90 0 0 la_oenb[58]
port 501 nsew signal input
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1120 90 0 0 la_oenb[59]
port 502 nsew signal input
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1120 90 0 0 la_oenb[5]
port 503 nsew signal input
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1120 90 0 0 la_oenb[60]
port 504 nsew signal input
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1120 90 0 0 la_oenb[61]
port 505 nsew signal input
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1120 90 0 0 la_oenb[62]
port 506 nsew signal input
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1120 90 0 0 la_oenb[63]
port 507 nsew signal input
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1120 90 0 0 la_oenb[64]
port 508 nsew signal input
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1120 90 0 0 la_oenb[65]
port 509 nsew signal input
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1120 90 0 0 la_oenb[66]
port 510 nsew signal input
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1120 90 0 0 la_oenb[67]
port 511 nsew signal input
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1120 90 0 0 la_oenb[68]
port 512 nsew signal input
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1120 90 0 0 la_oenb[69]
port 513 nsew signal input
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1120 90 0 0 la_oenb[6]
port 514 nsew signal input
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1120 90 0 0 la_oenb[70]
port 515 nsew signal input
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1120 90 0 0 la_oenb[71]
port 516 nsew signal input
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1120 90 0 0 la_oenb[72]
port 517 nsew signal input
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1120 90 0 0 la_oenb[73]
port 518 nsew signal input
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1120 90 0 0 la_oenb[74]
port 519 nsew signal input
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1120 90 0 0 la_oenb[75]
port 520 nsew signal input
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1120 90 0 0 la_oenb[76]
port 521 nsew signal input
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1120 90 0 0 la_oenb[77]
port 522 nsew signal input
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1120 90 0 0 la_oenb[78]
port 523 nsew signal input
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1120 90 0 0 la_oenb[79]
port 524 nsew signal input
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1120 90 0 0 la_oenb[7]
port 525 nsew signal input
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1120 90 0 0 la_oenb[80]
port 526 nsew signal input
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1120 90 0 0 la_oenb[81]
port 527 nsew signal input
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1120 90 0 0 la_oenb[82]
port 528 nsew signal input
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1120 90 0 0 la_oenb[83]
port 529 nsew signal input
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1120 90 0 0 la_oenb[84]
port 530 nsew signal input
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1120 90 0 0 la_oenb[85]
port 531 nsew signal input
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1120 90 0 0 la_oenb[86]
port 532 nsew signal input
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1120 90 0 0 la_oenb[87]
port 533 nsew signal input
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1120 90 0 0 la_oenb[88]
port 534 nsew signal input
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1120 90 0 0 la_oenb[89]
port 535 nsew signal input
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1120 90 0 0 la_oenb[8]
port 536 nsew signal input
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1120 90 0 0 la_oenb[90]
port 537 nsew signal input
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1120 90 0 0 la_oenb[91]
port 538 nsew signal input
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1120 90 0 0 la_oenb[92]
port 539 nsew signal input
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1120 90 0 0 la_oenb[93]
port 540 nsew signal input
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1120 90 0 0 la_oenb[94]
port 541 nsew signal input
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1120 90 0 0 la_oenb[95]
port 542 nsew signal input
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1120 90 0 0 la_oenb[96]
port 543 nsew signal input
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1120 90 0 0 la_oenb[97]
port 544 nsew signal input
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1120 90 0 0 la_oenb[98]
port 545 nsew signal input
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1120 90 0 0 la_oenb[99]
port 546 nsew signal input
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1120 90 0 0 la_oenb[9]
port 547 nsew signal input
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1120 90 0 0 user_clock2
port 548 nsew signal input
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1120 90 0 0 user_irq[0]
port 549 nsew signal tristate
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1120 90 0 0 user_irq[1]
port 550 nsew signal tristate
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1120 90 0 0 user_irq[2]
port 551 nsew signal tristate
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1120 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1120 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1120 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1120 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1120 0 0 0 vdda1
port 556 nsew signal bidirectional
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1120 0 0 0 vdda1
port 557 nsew signal bidirectional
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1120 0 0 0 vdda1
port 558 nsew signal bidirectional
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1120 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1120 0 0 0 vdda2
port 560 nsew signal bidirectional
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1120 0 0 0 vdda2
port 561 nsew signal bidirectional
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 1920 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 1920 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1120 0 0 0 vssa1
port 564 nsew signal bidirectional
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1120 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1120 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1120 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1120 0 0 0 vssd1
port 568 nsew signal bidirectional
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1120 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1120 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1120 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal2 s 524 -800 636 480 0 FreeSans 1120 90 0 0 wb_clk_i
port 572 nsew signal input
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1120 90 0 0 wb_rst_i
port 573 nsew signal input
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1120 90 0 0 wbs_ack_o
port 574 nsew signal tristate
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1120 90 0 0 wbs_adr_i[0]
port 575 nsew signal input
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1120 90 0 0 wbs_adr_i[10]
port 576 nsew signal input
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1120 90 0 0 wbs_adr_i[11]
port 577 nsew signal input
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1120 90 0 0 wbs_adr_i[12]
port 578 nsew signal input
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1120 90 0 0 wbs_adr_i[13]
port 579 nsew signal input
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1120 90 0 0 wbs_adr_i[14]
port 580 nsew signal input
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1120 90 0 0 wbs_adr_i[15]
port 581 nsew signal input
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1120 90 0 0 wbs_adr_i[16]
port 582 nsew signal input
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1120 90 0 0 wbs_adr_i[17]
port 583 nsew signal input
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1120 90 0 0 wbs_adr_i[18]
port 584 nsew signal input
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1120 90 0 0 wbs_adr_i[19]
port 585 nsew signal input
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1120 90 0 0 wbs_adr_i[1]
port 586 nsew signal input
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1120 90 0 0 wbs_adr_i[20]
port 587 nsew signal input
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1120 90 0 0 wbs_adr_i[21]
port 588 nsew signal input
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1120 90 0 0 wbs_adr_i[22]
port 589 nsew signal input
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1120 90 0 0 wbs_adr_i[23]
port 590 nsew signal input
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1120 90 0 0 wbs_adr_i[24]
port 591 nsew signal input
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1120 90 0 0 wbs_adr_i[25]
port 592 nsew signal input
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1120 90 0 0 wbs_adr_i[26]
port 593 nsew signal input
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1120 90 0 0 wbs_adr_i[27]
port 594 nsew signal input
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1120 90 0 0 wbs_adr_i[28]
port 595 nsew signal input
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1120 90 0 0 wbs_adr_i[29]
port 596 nsew signal input
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1120 90 0 0 wbs_adr_i[2]
port 597 nsew signal input
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1120 90 0 0 wbs_adr_i[30]
port 598 nsew signal input
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1120 90 0 0 wbs_adr_i[31]
port 599 nsew signal input
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1120 90 0 0 wbs_adr_i[3]
port 600 nsew signal input
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1120 90 0 0 wbs_adr_i[4]
port 601 nsew signal input
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1120 90 0 0 wbs_adr_i[5]
port 602 nsew signal input
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1120 90 0 0 wbs_adr_i[6]
port 603 nsew signal input
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1120 90 0 0 wbs_adr_i[7]
port 604 nsew signal input
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1120 90 0 0 wbs_adr_i[8]
port 605 nsew signal input
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1120 90 0 0 wbs_adr_i[9]
port 606 nsew signal input
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1120 90 0 0 wbs_cyc_i
port 607 nsew signal input
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1120 90 0 0 wbs_dat_i[0]
port 608 nsew signal input
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1120 90 0 0 wbs_dat_i[10]
port 609 nsew signal input
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1120 90 0 0 wbs_dat_i[11]
port 610 nsew signal input
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1120 90 0 0 wbs_dat_i[12]
port 611 nsew signal input
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1120 90 0 0 wbs_dat_i[13]
port 612 nsew signal input
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1120 90 0 0 wbs_dat_i[14]
port 613 nsew signal input
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1120 90 0 0 wbs_dat_i[15]
port 614 nsew signal input
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1120 90 0 0 wbs_dat_i[16]
port 615 nsew signal input
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1120 90 0 0 wbs_dat_i[17]
port 616 nsew signal input
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1120 90 0 0 wbs_dat_i[18]
port 617 nsew signal input
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1120 90 0 0 wbs_dat_i[19]
port 618 nsew signal input
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1120 90 0 0 wbs_dat_i[1]
port 619 nsew signal input
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1120 90 0 0 wbs_dat_i[20]
port 620 nsew signal input
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1120 90 0 0 wbs_dat_i[21]
port 621 nsew signal input
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1120 90 0 0 wbs_dat_i[22]
port 622 nsew signal input
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1120 90 0 0 wbs_dat_i[23]
port 623 nsew signal input
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1120 90 0 0 wbs_dat_i[24]
port 624 nsew signal input
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1120 90 0 0 wbs_dat_i[25]
port 625 nsew signal input
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1120 90 0 0 wbs_dat_i[26]
port 626 nsew signal input
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1120 90 0 0 wbs_dat_i[27]
port 627 nsew signal input
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1120 90 0 0 wbs_dat_i[28]
port 628 nsew signal input
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1120 90 0 0 wbs_dat_i[29]
port 629 nsew signal input
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1120 90 0 0 wbs_dat_i[2]
port 630 nsew signal input
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1120 90 0 0 wbs_dat_i[30]
port 631 nsew signal input
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1120 90 0 0 wbs_dat_i[31]
port 632 nsew signal input
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1120 90 0 0 wbs_dat_i[3]
port 633 nsew signal input
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1120 90 0 0 wbs_dat_i[4]
port 634 nsew signal input
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1120 90 0 0 wbs_dat_i[5]
port 635 nsew signal input
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1120 90 0 0 wbs_dat_i[6]
port 636 nsew signal input
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1120 90 0 0 wbs_dat_i[7]
port 637 nsew signal input
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1120 90 0 0 wbs_dat_i[8]
port 638 nsew signal input
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1120 90 0 0 wbs_dat_i[9]
port 639 nsew signal input
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1120 90 0 0 wbs_dat_o[0]
port 640 nsew signal tristate
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1120 90 0 0 wbs_dat_o[10]
port 641 nsew signal tristate
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1120 90 0 0 wbs_dat_o[11]
port 642 nsew signal tristate
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1120 90 0 0 wbs_dat_o[12]
port 643 nsew signal tristate
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1120 90 0 0 wbs_dat_o[13]
port 644 nsew signal tristate
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1120 90 0 0 wbs_dat_o[14]
port 645 nsew signal tristate
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1120 90 0 0 wbs_dat_o[15]
port 646 nsew signal tristate
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1120 90 0 0 wbs_dat_o[16]
port 647 nsew signal tristate
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1120 90 0 0 wbs_dat_o[17]
port 648 nsew signal tristate
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1120 90 0 0 wbs_dat_o[18]
port 649 nsew signal tristate
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1120 90 0 0 wbs_dat_o[19]
port 650 nsew signal tristate
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1120 90 0 0 wbs_dat_o[1]
port 651 nsew signal tristate
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1120 90 0 0 wbs_dat_o[20]
port 652 nsew signal tristate
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1120 90 0 0 wbs_dat_o[21]
port 653 nsew signal tristate
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1120 90 0 0 wbs_dat_o[22]
port 654 nsew signal tristate
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1120 90 0 0 wbs_dat_o[23]
port 655 nsew signal tristate
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1120 90 0 0 wbs_dat_o[24]
port 656 nsew signal tristate
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1120 90 0 0 wbs_dat_o[25]
port 657 nsew signal tristate
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1120 90 0 0 wbs_dat_o[26]
port 658 nsew signal tristate
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1120 90 0 0 wbs_dat_o[27]
port 659 nsew signal tristate
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1120 90 0 0 wbs_dat_o[28]
port 660 nsew signal tristate
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1120 90 0 0 wbs_dat_o[29]
port 661 nsew signal tristate
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1120 90 0 0 wbs_dat_o[2]
port 662 nsew signal tristate
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1120 90 0 0 wbs_dat_o[30]
port 663 nsew signal tristate
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1120 90 0 0 wbs_dat_o[31]
port 664 nsew signal tristate
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1120 90 0 0 wbs_dat_o[3]
port 665 nsew signal tristate
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1120 90 0 0 wbs_dat_o[4]
port 666 nsew signal tristate
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1120 90 0 0 wbs_dat_o[5]
port 667 nsew signal tristate
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1120 90 0 0 wbs_dat_o[6]
port 668 nsew signal tristate
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1120 90 0 0 wbs_dat_o[7]
port 669 nsew signal tristate
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1120 90 0 0 wbs_dat_o[8]
port 670 nsew signal tristate
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1120 90 0 0 wbs_dat_o[9]
port 671 nsew signal tristate
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1120 90 0 0 wbs_sel_i[0]
port 672 nsew signal input
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1120 90 0 0 wbs_sel_i[1]
port 673 nsew signal input
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1120 90 0 0 wbs_sel_i[2]
port 674 nsew signal input
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1120 90 0 0 wbs_sel_i[3]
port 675 nsew signal input
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1120 90 0 0 wbs_stb_i
port 676 nsew signal input
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1120 90 0 0 wbs_we_i
port 677 nsew signal input
rlabel metal5 564246 213496 568826 217492 1 gnd
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
