magic
tech sky130A
magscale 1 2
timestamp 1672355014
<< error_p >>
rect -30 130 30 136
rect -30 97 -18 130
rect -30 96 18 97
rect -30 90 30 96
rect 34 -49 36 50
rect -34 -50 36 -49
rect -30 -96 30 -90
rect -30 -130 -18 -96
rect -30 -136 30 -130
<< nwell >>
rect -230 -268 230 268
<< pmoslvt >>
rect -34 -50 34 50
<< pdiff >>
rect -92 38 -34 50
rect -92 -38 -80 38
rect -46 -38 -34 38
rect -92 -50 -34 -38
rect 34 38 92 50
rect 34 -38 46 38
rect 80 -38 92 38
rect 34 -50 92 -38
<< pdiffc >>
rect -80 -38 -46 38
rect 46 -38 80 38
<< nsubdiff >>
rect -194 198 -98 232
rect 98 198 194 232
rect -194 136 -160 198
rect 160 136 194 198
rect -194 -198 -160 -136
rect 160 -198 194 -136
rect -194 -232 -98 -198
rect 98 -232 194 -198
<< nsubdiffcont >>
rect -98 198 98 232
rect -194 -136 -160 136
rect 160 -136 194 136
rect -98 -232 98 -198
<< poly >>
rect -34 130 34 146
rect -34 96 -18 130
rect 18 96 34 130
rect -34 50 34 96
rect -34 -96 34 -50
rect -34 -130 -18 -96
rect 18 -130 34 -96
rect -34 -146 34 -130
<< polycont >>
rect -18 96 18 130
rect -18 -130 18 -96
<< locali >>
rect -194 198 -98 232
rect 98 198 194 232
rect -194 136 -160 198
rect 160 136 194 198
rect -34 96 -18 130
rect 18 96 34 130
rect -80 38 -46 54
rect -80 -54 -46 -38
rect 46 38 80 54
rect 46 -54 80 -38
rect -34 -130 -18 -96
rect 18 -130 34 -96
rect -194 -198 -160 -136
rect 160 -198 194 -136
rect -194 -232 -98 -198
rect 98 -232 194 -198
<< viali >>
rect -18 96 18 130
rect -80 -38 -46 38
rect 46 -38 80 38
rect -18 -130 18 -96
<< metal1 >>
rect -30 130 30 136
rect -30 96 -18 130
rect 18 96 30 130
rect -30 90 30 96
rect -86 38 -40 50
rect -86 -38 -80 38
rect -46 -38 -40 38
rect -86 -50 -40 -38
rect 40 38 86 50
rect 40 -38 46 38
rect 80 -38 86 38
rect 40 -50 86 -38
rect -30 -96 30 -90
rect -30 -130 -18 -96
rect 18 -130 30 -96
rect -30 -136 30 -130
<< properties >>
string FIXED_BBOX -178 -216 178 216
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 0.5 l 0.35 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
