magic
tech sky130A
magscale 1 2
timestamp 1672466235
<< locali >>
rect 18631 -14326 18677 -13625
rect 18631 -14372 24739 -14326
rect 18946 -34170 21745 -34124
rect 21791 -34170 25561 -34124
rect 19385 -38985 19475 -38875
rect 19105 -38991 19475 -38985
rect 19105 -39069 19111 -38991
rect 19189 -39069 19475 -38991
rect 19105 -39075 19475 -39069
rect 19385 -41125 19475 -39075
rect 21015 -41125 21105 -38805
rect 19385 -41215 21105 -41125
<< viali >>
rect 24739 -14372 24785 -14326
rect 21745 -34170 21791 -34124
rect 19111 -39069 19189 -38991
<< metal1 >>
rect 17860 -14314 19206 -13638
rect 21080 -14110 21775 -13640
rect 22245 -14110 22251 -13640
rect 21080 -14250 21550 -14110
rect 24727 -14326 24797 -14320
rect 24727 -14378 24733 -14326
rect 24791 -14378 24797 -14326
rect 24733 -14384 24791 -14378
rect 21449 -33209 21631 -33203
rect 21631 -33391 25481 -33209
rect 21449 -33397 21631 -33391
rect 18564 -34070 18570 -33870
rect 18770 -34070 19620 -33870
rect 20970 -33930 21460 -33900
rect 25299 -33920 25481 -33391
rect 20970 -34050 23230 -33930
rect 20975 -34080 23230 -34050
rect 24990 -34061 25481 -33920
rect 24990 -34070 25480 -34061
rect 21733 -34124 21803 -34118
rect 21733 -34176 21739 -34124
rect 21797 -34176 21803 -34124
rect 21739 -34182 21797 -34176
rect 22015 -34425 22165 -34080
rect 26205 -34425 26355 -34419
rect 22015 -34575 26205 -34425
rect 26205 -34581 26355 -34575
rect 21184 -37620 21190 -37460
rect 21350 -37620 21356 -37460
rect 19330 -37750 19460 -37744
rect 19460 -37880 20325 -37750
rect 19330 -37886 19460 -37880
rect 20195 -38225 20325 -37880
rect 20195 -38355 20905 -38225
rect 19600 -38940 19700 -38450
rect 20775 -38935 20905 -38355
rect 21190 -38970 21350 -37620
rect 20213 -38980 20307 -38978
rect 20710 -38980 20800 -38970
rect 19500 -38985 19590 -38980
rect 19099 -38991 19590 -38985
rect 19099 -39069 19111 -38991
rect 19189 -39069 19590 -38991
rect 19099 -39075 19590 -39069
rect 19500 -40990 19590 -39075
rect 19710 -39070 20800 -38980
rect 19710 -40990 19800 -39070
rect 20213 -46463 20307 -39070
rect 20710 -40980 20800 -39070
rect 20910 -39130 21350 -38970
rect 20910 -40980 21000 -39130
rect 21617 -46463 21623 -46462
rect 20213 -46557 21623 -46463
rect 21718 -46557 21724 -46462
<< via1 >>
rect 21775 -14110 22245 -13640
rect 24733 -14372 24739 -14326
rect 24739 -14372 24785 -14326
rect 24785 -14372 24791 -14326
rect 24733 -14378 24791 -14372
rect 21449 -33391 21631 -33209
rect 18570 -34070 18770 -33870
rect 21739 -34170 21745 -34124
rect 21745 -34170 21791 -34124
rect 21791 -34170 21797 -34124
rect 21739 -34176 21797 -34170
rect 26205 -34575 26355 -34425
rect 21190 -37620 21350 -37460
rect 19330 -37880 19460 -37750
rect 21623 -46557 21718 -46462
<< metal2 >>
rect 21775 -13640 22245 -13631
rect 21775 -14119 22245 -14110
rect 24732 -14322 24792 -14313
rect 24727 -14378 24732 -14326
rect 24792 -14378 24797 -14326
rect 24732 -14391 24792 -14382
rect 21454 -33209 21626 -33205
rect 21443 -33391 21449 -33209
rect 21631 -33391 21637 -33209
rect 21454 -33395 21626 -33391
rect 18570 -33870 18770 -33861
rect 18570 -34079 18770 -34070
rect 21738 -34120 21798 -34111
rect 21733 -34176 21738 -34124
rect 21798 -34176 21803 -34124
rect 21738 -34189 21798 -34180
rect 26205 -34425 26355 -34416
rect 26199 -34575 26205 -34425
rect 26355 -34575 26361 -34425
rect 26205 -34584 26355 -34575
rect 21190 -37460 21350 -37454
rect 21186 -37615 21190 -37465
rect 21350 -37615 21354 -37465
rect 21190 -37626 21350 -37620
rect 19335 -37750 19455 -37746
rect 19324 -37880 19330 -37750
rect 19460 -37880 19466 -37750
rect 19335 -37884 19455 -37880
rect 21623 -46462 21718 -46456
rect 21614 -46557 21623 -46462
rect 21718 -46557 21727 -46462
rect 21623 -46563 21718 -46557
<< via2 >>
rect 21775 -14110 22245 -13640
rect 24732 -14326 24792 -14322
rect 24732 -14378 24733 -14326
rect 24733 -14378 24791 -14326
rect 24791 -14378 24792 -14326
rect 24732 -14382 24792 -14378
rect 21454 -33386 21626 -33214
rect 18570 -34070 18770 -33870
rect 21738 -34124 21798 -34120
rect 21738 -34176 21739 -34124
rect 21739 -34176 21797 -34124
rect 21797 -34176 21798 -34124
rect 21738 -34180 21798 -34176
rect 26205 -34575 26355 -34425
rect 21195 -37615 21345 -37465
rect 19335 -37875 19455 -37755
rect 21623 -46557 21718 -46462
<< metal3 >>
rect 21770 -13640 22250 -13635
rect 21770 -13645 21775 -13640
rect 22245 -13645 22250 -13640
rect 21770 -14121 22250 -14115
rect 24727 -14322 24797 -14317
rect 24727 -14382 24732 -14322
rect 24792 -14382 24797 -14322
rect 24727 -14387 24797 -14382
rect 24732 -14840 24792 -14387
rect 24670 -32960 24850 -14840
rect 24600 -33060 24850 -32960
rect 21450 -33209 21630 -33204
rect 21449 -33210 21631 -33209
rect 21449 -33390 21450 -33210
rect 21630 -33390 21631 -33210
rect 24600 -33360 24840 -33060
rect 21449 -33391 21631 -33390
rect 21450 -33396 21630 -33391
rect 22040 -33528 24840 -33360
rect 18190 -33600 24840 -33528
rect 18190 -33768 22280 -33600
rect 18190 -35222 18430 -33768
rect 18559 -34075 18565 -33865
rect 18765 -33870 18775 -33865
rect 18770 -34070 18775 -33870
rect 18765 -34075 18775 -34070
rect 21738 -34115 21798 -33768
rect 22040 -33804 22280 -33768
rect 21733 -34120 21803 -34115
rect 21733 -34180 21738 -34120
rect 21798 -34180 21803 -34120
rect 21733 -34185 21803 -34180
rect 21738 -34220 21798 -34185
rect 26200 -34425 26360 -34420
rect 26200 -34575 26205 -34425
rect 26355 -34575 26360 -34425
rect 26200 -34580 26360 -34575
rect 26205 -35125 26355 -34580
rect 20870 -37465 21350 -37460
rect 20870 -37615 21195 -37465
rect 21345 -37615 21350 -37465
rect 20870 -37620 21350 -37615
rect 19331 -37750 19459 -37745
rect 19330 -37751 19460 -37750
rect 19330 -37879 19331 -37751
rect 19459 -37879 19460 -37751
rect 19330 -37880 19460 -37879
rect 19331 -37885 19459 -37880
rect 21618 -46462 21628 -46457
rect 21618 -46557 21623 -46462
rect 21618 -46562 21628 -46557
rect 21723 -46562 21729 -46457
<< via3 >>
rect 21770 -14110 21775 -13645
rect 21775 -14110 22245 -13645
rect 22245 -14110 22250 -13645
rect 21770 -14115 22250 -14110
rect 21450 -33214 21630 -33210
rect 21450 -33386 21454 -33214
rect 21454 -33386 21626 -33214
rect 21626 -33386 21630 -33214
rect 21450 -33390 21630 -33386
rect 18565 -33870 18765 -33865
rect 18565 -34070 18570 -33870
rect 18570 -34070 18765 -33870
rect 18565 -34075 18765 -34070
rect 19331 -37755 19459 -37751
rect 19331 -37875 19335 -37755
rect 19335 -37875 19455 -37755
rect 19455 -37875 19459 -37755
rect 19331 -37879 19459 -37875
rect 21628 -46462 21723 -46457
rect 21628 -46557 21718 -46462
rect 21718 -46557 21723 -46462
rect 21628 -46562 21723 -46557
<< metal4 >>
rect 21769 -13645 22251 -13644
rect 21769 -14115 21770 -13645
rect 22250 -14115 22251 -13645
rect 21769 -14116 22251 -14115
rect 21775 -15495 22245 -14116
rect 21449 -33210 21631 -32829
rect 21449 -33390 21450 -33210
rect 21630 -33390 21631 -33210
rect 21449 -33391 21631 -33390
rect 18564 -33865 18766 -33864
rect 18564 -34075 18565 -33865
rect 18765 -34075 18766 -33865
rect 18564 -34076 18766 -34075
rect 18565 -35040 18765 -34076
rect 19330 -37751 19460 -37420
rect 19330 -37879 19331 -37751
rect 19459 -37879 19460 -37751
rect 19330 -37880 19460 -37879
rect 21627 -46457 21724 -46456
rect 21627 -46562 21628 -46457
rect 21723 -46461 21724 -46457
rect 21723 -46556 22267 -46461
rect 21723 -46562 21724 -46556
rect 21627 -46563 21724 -46562
use sky130_fd_pr__cap_mim_m3_1_4BCNTW  XC4
timestamp 1672466235
transform 1 0 24186 0 1 -41080
box -2186 -6320 2186 6320
use sky130_fd_pr__cap_mim_m3_1_NUYDZ7  XC27
timestamp 1672466235
transform 1 0 21686 0 1 -24020
box -3086 -9180 3086 9180
use sky130_fd_pr__res_xhigh_po_2p85_QPY2BD  XR7
timestamp 1672466235
transform 0 1 20148 -1 0 -13949
box -450 -1548 450 1548
use sky130_fd_pr__res_xhigh_po_0p69_LVNRZ4  XR23
timestamp 1672466235
transform 0 1 20288 -1 0 -33965
box -234 -1288 234 1288
use sky130_fd_pr__cap_mim_m3_1_TE3E2R  sky130_fd_pr__cap_mim_m3_1_TE3E2R_0
timestamp 1672466235
transform 1 0 19574 0 1 -36072
box -1587 -1441 1587 1441
use sky130_fd_pr__pfet_01v8_lvt_8R53B2  sky130_fd_pr__pfet_01v8_lvt_8R53B2_0
timestamp 1672466235
transform 1 0 19649 0 1 -39981
box -247 -1219 247 1219
use sky130_fd_pr__pfet_01v8_lvt_8R53B2  sky130_fd_pr__pfet_01v8_lvt_X3MKZ5_0
timestamp 1672466235
transform 1 0 20849 0 1 -39981
box -247 -1219 247 1219
use sky130_fd_pr__res_xhigh_po_0p35_4XRDQ9  sky130_fd_pr__res_xhigh_po_0p35_4XRDQ9_0
timestamp 1672466235
transform 0 1 24130 -1 0 -34009
box -201 -1498 201 1498
<< labels >>
rlabel metal1 18018 -14164 18352 -13744 1 input
port 1 n
rlabel metal1 21236 -39054 21264 -38898 1 gnd
port 4 n
rlabel metal1 19232 -39058 19270 -39030 1 vcc
port 0 n
rlabel metal1 19610 -38612 19688 -38568 1 pb
port 3 n
rlabel metal1 20226 -39058 20304 -39014 1 out
port 2 n
<< end >>
