magic
tech sky130A
magscale 1 2
timestamp 1672366615
<< locali >>
rect -4360 5304 11420 5310
rect -4360 5216 256 5304
rect 344 5216 11420 5304
rect -4360 5210 11420 5216
rect -20 4310 80 5210
rect -4340 4210 11390 4310
rect -40 3050 60 4210
rect -2560 2950 60 3050
rect 1169 2100 1210 2960
rect 1029 2059 1210 2100
rect 1029 1750 1070 2059
rect 1375 1959 12785 1965
rect 1375 1921 12741 1959
rect 12779 1921 12785 1959
rect 1375 1915 12785 1921
rect -1890 1709 1070 1750
rect -1890 1591 -1849 1709
rect -2480 1550 -1190 1591
rect -1890 457 -1850 1550
rect 1029 871 1070 1709
rect -1890 423 -1887 457
rect -1853 423 -1850 457
rect -1890 270 -1850 423
rect -2490 230 -1230 270
rect -1890 190 -1850 230
<< viali >>
rect 256 5216 344 5304
rect 1325 1915 1375 1965
rect 12741 1921 12779 1959
rect 1029 830 1070 871
rect -1887 423 -1853 457
rect -1890 150 -1850 190
<< metal1 >>
rect -4180 5500 11240 6080
rect -4180 5110 -3590 5500
rect -2330 5160 -880 5500
rect 250 5304 350 5500
rect 250 5216 256 5304
rect 344 5216 350 5304
rect 250 5204 350 5216
rect 1670 5160 10760 5500
rect -2580 5100 -580 5160
rect -4315 4635 -4225 5085
rect -3540 5010 -2620 5080
rect -4180 4900 -3590 4990
rect -2580 4900 -580 4990
rect -540 4980 1170 5110
rect 1220 5100 11220 5160
rect 11270 5010 11300 5080
rect -3895 4635 -3805 4900
rect -4315 4545 -3805 4635
rect -3895 4200 -3805 4545
rect -2580 4200 -2490 4900
rect -680 4200 -590 4900
rect -4170 4110 -3580 4200
rect -2590 4110 -590 4200
rect 1210 4700 11220 4990
rect 1210 4400 1500 4700
rect 10905 4400 11195 4700
rect 1210 4110 11220 4400
rect -4295 3565 -4225 4085
rect -3540 4010 -2630 4080
rect -4180 3920 -3580 3990
rect -3905 3565 -3835 3920
rect -2580 3900 -580 3990
rect -540 3980 1170 4110
rect 11270 4010 11300 4080
rect -4295 3495 -3735 3565
rect -3805 3160 -3735 3495
rect -1575 3455 -1485 3900
rect 1220 3540 11200 4000
rect 1220 3520 1680 3540
rect -1865 3365 -1485 3455
rect -3860 2460 -3680 3160
rect -2690 2860 -2310 2910
rect -2485 2295 -2415 2815
rect -2705 2225 -2415 2295
rect -2290 2805 -2220 2810
rect -1865 2805 -1775 3365
rect -1400 2860 -1020 2910
rect -2290 2735 -1415 2805
rect -2290 2230 -2220 2735
rect -2705 1710 -2635 2225
rect -1485 2215 -1415 2735
rect -1295 2285 -1225 2815
rect 1210 2655 1720 2940
rect 615 2585 1720 2655
rect -1295 2215 -975 2285
rect -1045 1825 -975 2215
rect 615 1825 685 2585
rect 1210 2350 1720 2585
rect 3740 2690 4250 2910
rect 10740 2870 11200 3540
rect 3740 2580 4625 2690
rect 4735 2580 4741 2690
rect 3740 2320 4250 2580
rect 7694 2410 7700 2870
rect 8160 2410 13580 2870
rect 1319 1965 1381 1977
rect 1105 1915 1325 1965
rect 1375 1915 1381 1965
rect -1045 1755 695 1825
rect -2705 1670 -2030 1710
rect -2705 1400 -2635 1670
rect -2070 1490 -2030 1670
rect -2400 1450 -1310 1490
rect -2705 1390 -2410 1400
rect -2710 1330 -2410 1390
rect -3830 140 -3430 390
rect -2710 370 -2670 1330
rect -2480 420 -2410 1330
rect -2290 460 -2250 1410
rect -1893 460 -1847 463
rect -1450 460 -1410 1410
rect -1045 1400 -975 1755
rect 625 1555 695 1755
rect 1105 1555 1155 1915
rect 1319 1903 1381 1915
rect 10740 1760 11200 2410
rect 12729 1959 13255 1965
rect 12729 1921 12741 1959
rect 12779 1921 13255 1959
rect 12729 1915 13255 1921
rect 625 1485 1175 1555
rect -2300 457 -1410 460
rect -2300 423 -1887 457
rect -1853 423 -1410 457
rect -2300 420 -1410 423
rect -1300 1330 -975 1400
rect -1300 420 -1230 1330
rect 1105 1185 1175 1485
rect 1220 1300 13010 1760
rect 13040 1230 13090 1290
rect 13205 1230 13255 1915
rect 1210 1140 13000 1200
rect 13040 1180 13255 1230
rect 1410 1130 13000 1140
rect 1410 1000 12800 1130
rect 1210 990 12800 1000
rect 1017 871 1082 877
rect 1210 871 13040 990
rect 1017 830 1029 871
rect 1070 830 13040 871
rect 1017 824 1082 830
rect -1893 417 -1847 420
rect -2710 330 -1310 370
rect -1896 190 -1844 202
rect 1210 190 13040 830
rect -1896 150 -1890 190
rect -1850 150 13040 190
rect -1896 140 13040 150
rect -3830 -50 1590 140
rect -3500 -60 1590 -50
<< via1 >>
rect 4625 2580 4735 2690
rect 7700 2410 8160 2870
<< metal2 >>
rect 7700 2870 8160 2876
rect 4625 2690 4735 2696
rect 4616 2580 4625 2690
rect 4735 2580 4744 2690
rect 4625 2574 4735 2580
rect 7691 2410 7700 2870
rect 8160 2410 8169 2870
rect 7700 2404 8160 2410
<< via2 >>
rect 4625 2580 4735 2690
rect 7700 2410 8160 2870
<< metal3 >>
rect 4620 2690 4740 2695
rect 4620 2580 4625 2690
rect 4735 2580 5375 2690
rect 4620 2575 4740 2580
rect 7689 2405 7695 2875
rect 8155 2870 8165 2875
rect 8160 2410 8165 2870
rect 8155 2405 8165 2410
<< via3 >>
rect 7695 2870 8155 2875
rect 7695 2410 7700 2870
rect 7700 2410 8155 2870
rect 7695 2405 8155 2410
<< metal4 >>
rect 7694 2875 8156 2876
rect 7694 2870 7695 2875
rect 6230 2410 7695 2870
rect 7694 2405 7695 2410
rect 8155 2405 8156 2875
rect 7694 2404 8156 2405
use sky130_fd_pr__cap_mim_m3_1_KYM84V  XC6
timestamp 1672354625
transform -1 0 6016 0 -1 2600
box -886 -740 886 740
use sky130_fd_pr__pfet_01v8_lvt_XP5BXZ  XM53
timestamp 1672366615
transform 0 -1 -3881 1 0 5050
box -247 -519 247 519
use sky130_fd_pr__pfet_01v8_lvt_XP5BXZ  XM54
timestamp 1672366615
transform 1 0 -2350 0 1 2519
box -247 -519 247 519
use sky130_fd_pr__pfet_01v8_lvt_X3MKZ5  XM56
timestamp 1672354625
transform 0 -1 -1581 1 0 5046
box -246 -1219 246 1219
use sky130_fd_pr__nfet_01v8_lvt_MYKW3H  XM57
timestamp 1672354625
transform 0 1 7110 -1 0 1246
box -246 -6110 246 6110
use sky130_fd_pr__pfet_01v8_lvt_X3MKZ5  XM59
timestamp 1672354625
transform 0 -1 -1581 1 0 4046
box -246 -1219 246 1219
use sky130_fd_pr__nfet_01v8_lvt_8TEW3F  XM60
timestamp 1672354625
transform 1 0 -2354 0 1 910
box -246 -710 246 710
use sky130_fd_pr__nfet_01v8_lvt_8TEW3F  XM61
timestamp 1672354625
transform 1 0 -1354 0 1 910
box -246 -710 246 710
use sky130_fd_pr__pfet_01v8_lvt_X3MVBA  XM62
timestamp 1672354625
transform 0 1 6219 -1 0 5046
box -246 -5219 246 5219
use sky130_fd_pr__pfet_01v8_lvt_X3MVBA  XM63
timestamp 1672354625
transform 0 1 6219 -1 0 4046
box -246 -5219 246 5219
use sky130_fd_pr__res_xhigh_po_0p69_FR2N8V  XR17
timestamp 1672354625
transform 1 0 -3765 0 1 1438
box -234 -1638 234 1638
use sky130_fd_pr__res_high_po_2p85_HV4VUF  XR18
timestamp 1672354625
transform 0 -1 2738 1 0 2621
box -450 -1598 450 1598
use sky130_fd_pr__pfet_01v8_lvt_XP5BXZ  sky130_fd_pr__pfet_01v8_lvt_XP5BXZ_0
timestamp 1672366615
transform 0 -1 -3881 1 0 4050
box -247 -519 247 519
use sky130_fd_pr__pfet_01v8_lvt_XP5BXZ  sky130_fd_pr__pfet_01v8_lvt_XP5BXZ_1
timestamp 1672366615
transform 1 0 -1350 0 1 2519
box -247 -519 247 519
<< labels >>
rlabel metal1 -1200 5690 -1090 5840 1 vcc
port 0 n
rlabel metal1 -2670 2880 -2640 2900 1 inv
port 1 n
rlabel metal1 -1080 2870 -1050 2890 1 noninv
port 2 n
rlabel metal1 12440 2630 12470 2650 1 output
port 3 n
rlabel metal1 4864 332 4938 422 1 gnd
port 4 n
<< end >>
