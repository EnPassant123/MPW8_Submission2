magic
tech sky130A
timestamp 1672002055
<< metal3 >>
rect -2726 2566 -60 2580
rect -2726 74 -102 2566
rect -70 74 -60 2566
rect -2726 60 -60 74
rect 60 2566 2726 2580
rect 60 74 2684 2566
rect 2716 74 2726 2566
rect 60 60 2726 74
rect -2726 -74 -60 -60
rect -2726 -2566 -102 -74
rect -70 -2566 -60 -74
rect -2726 -2580 -60 -2566
rect 60 -74 2726 -60
rect 60 -2566 2684 -74
rect 2716 -2566 2726 -74
rect 60 -2580 2726 -2566
<< via3 >>
rect -102 74 -70 2566
rect 2684 74 2716 2566
rect -102 -2566 -70 -74
rect 2684 -2566 2716 -74
<< mimcap >>
rect -2706 2540 -226 2560
rect -2706 100 -2686 2540
rect -246 100 -226 2540
rect -2706 80 -226 100
rect 80 2540 2560 2560
rect 80 100 100 2540
rect 2540 100 2560 2540
rect 80 80 2560 100
rect -2706 -100 -226 -80
rect -2706 -2540 -2686 -100
rect -246 -2540 -226 -100
rect -2706 -2560 -226 -2540
rect 80 -100 2560 -80
rect 80 -2540 100 -100
rect 2540 -2540 2560 -100
rect 80 -2560 2560 -2540
<< mimcapcontact >>
rect -2686 100 -246 2540
rect 100 100 2540 2540
rect -2686 -2540 -246 -100
rect 100 -2540 2540 -100
<< metal4 >>
rect -1492 2540 -1440 2640
rect -112 2566 -60 2640
rect -246 100 -245 2540
rect -2686 99 -245 100
rect -1492 -99 -1440 99
rect -112 74 -102 2566
rect -70 74 -60 2566
rect 1294 2540 1346 2640
rect 2674 2566 2726 2640
rect 99 100 100 2540
rect 99 99 2540 100
rect -112 -74 -60 74
rect -2686 -100 -245 -99
rect -246 -2540 -245 -100
rect -1492 -2640 -1440 -2540
rect -112 -2566 -102 -74
rect -70 -2566 -60 -74
rect 1294 -99 1346 99
rect 2674 74 2684 2566
rect 2716 74 2726 2566
rect 2674 -74 2726 74
rect 99 -100 2540 -99
rect 99 -2540 100 -100
rect -112 -2640 -60 -2566
rect 1294 -2640 1346 -2540
rect 2674 -2566 2684 -74
rect 2716 -2566 2726 -74
rect 2674 -2640 2726 -2566
<< properties >>
string FIXED_BBOX 60 60 2580 2580
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 24.8 l 24.8 val 1.248k carea 2.00 cperi 0.19 nx 2 ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
