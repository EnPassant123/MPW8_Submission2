magic
tech sky130A
magscale 1 2
timestamp 1672362834
<< pwell >>
rect -201 -3598 201 3598
<< psubdiff >>
rect -165 3528 -69 3562
rect 69 3528 165 3562
rect -165 3466 -131 3528
rect 131 3466 165 3528
rect -165 -3528 -131 -3466
rect 131 -3528 165 -3466
rect -165 -3562 -69 -3528
rect 69 -3562 165 -3528
<< psubdiffcont >>
rect -69 3528 69 3562
rect -165 -3466 -131 3466
rect 131 -3466 165 3466
rect -69 -3562 69 -3528
<< xpolycontact >>
rect -35 3000 35 3432
rect -35 -3432 35 -3000
<< xpolyres >>
rect -35 -3000 35 3000
<< locali >>
rect -165 3528 -69 3562
rect 69 3528 165 3562
rect -165 3466 -131 3528
rect 131 3466 165 3528
rect -165 -3528 -131 -3466
rect 131 -3528 165 -3466
rect -165 -3562 -69 -3528
rect 69 -3562 165 -3528
<< viali >>
rect -19 3017 19 3414
rect -19 -3414 19 -3017
<< metal1 >>
rect -25 3414 25 3426
rect -25 3017 -19 3414
rect 19 3017 25 3414
rect -25 3005 25 3017
rect -25 -3017 25 -3005
rect -25 -3414 -19 -3017
rect 19 -3414 25 -3017
rect -25 -3426 25 -3414
<< res0p35 >>
rect -37 -3002 37 3002
<< properties >>
string FIXED_BBOX -148 -3545 148 3545
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 29.995 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 172.475k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
