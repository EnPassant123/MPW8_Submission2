magic
tech sky130A
magscale 1 2
timestamp 1672353341
<< error_p >>
rect -34 446 34 447
rect -50 -400 50 -399
<< nwell >>
rect -246 -618 246 618
<< pmoslvt >>
rect -50 -400 50 400
<< pdiff >>
rect -108 388 -50 400
rect -108 -388 -96 388
rect -62 -388 -50 388
rect -108 -400 -50 -388
rect 50 388 108 400
rect 50 -388 62 388
rect 96 -388 108 388
rect 50 -400 108 -388
<< pdiffc >>
rect -96 -388 -62 388
rect 62 -388 96 388
<< nsubdiff >>
rect -210 548 -114 582
rect 114 548 210 582
rect -210 486 -176 548
rect 176 486 210 548
rect -210 -548 -176 -486
rect 176 -548 210 -486
rect -210 -582 -114 -548
rect 114 -582 210 -548
<< nsubdiffcont >>
rect -114 548 114 582
rect -210 -486 -176 486
rect 176 -486 210 486
rect -114 -582 114 -548
<< poly >>
rect -50 480 50 496
rect -50 446 -34 480
rect 34 446 50 480
rect -50 400 50 446
rect -50 -446 50 -400
rect -50 -480 -34 -446
rect 34 -480 50 -446
rect -50 -496 50 -480
<< polycont >>
rect -34 446 34 480
rect -34 -480 34 -446
<< locali >>
rect -210 548 -114 582
rect 114 548 210 582
rect -210 486 -176 548
rect 176 486 210 548
rect -50 446 -34 480
rect 34 446 50 480
rect -96 388 -62 404
rect -96 -404 -62 -388
rect 62 388 96 404
rect 62 -404 96 -388
rect -50 -480 -34 -446
rect 34 -480 50 -446
rect -210 -548 -176 -486
rect 176 -548 210 -486
rect -210 -582 -114 -548
rect 114 -582 210 -548
<< viali >>
rect -34 446 34 480
rect -96 -388 -62 388
rect 62 -388 96 388
rect -34 -480 34 -446
<< metal1 >>
rect -46 480 46 486
rect -46 446 -34 480
rect 34 446 46 480
rect -46 440 46 446
rect -102 388 -56 400
rect -102 -388 -96 388
rect -62 -388 -56 388
rect -102 -400 -56 -388
rect 56 388 102 400
rect 56 -388 62 388
rect 96 -388 102 388
rect 56 -400 102 -388
rect -46 -446 46 -440
rect -46 -480 -34 -446
rect 34 -480 46 -446
rect -46 -486 46 -480
<< properties >>
string FIXED_BBOX -192 -566 192 566
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 4.0 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
