magic
tech sky130A
timestamp 1671518644
<< pwell >>
rect -100 -749 100 749
<< psubdiff >>
rect -82 714 -34 731
rect 34 714 82 731
rect -82 683 -65 714
rect 65 683 82 714
rect -82 -714 -65 -683
rect 65 -714 82 -683
rect -82 -731 -34 -714
rect 34 -731 82 -714
<< psubdiffcont >>
rect -34 714 34 731
rect -82 -683 -65 683
rect 65 -683 82 683
rect -34 -731 34 -714
<< xpolycontact >>
rect -17 450 17 666
rect -17 -666 17 -450
<< xpolyres >>
rect -17 -450 17 450
<< locali >>
rect -82 714 -34 731
rect 34 714 82 731
rect -82 683 -65 714
rect 65 683 82 714
rect -82 -714 -65 -683
rect 65 -714 82 -683
rect -82 -731 -34 -714
rect 34 -731 82 -714
<< viali >>
rect -9 458 9 657
rect -9 -657 9 -458
<< metal1 >>
rect -12 657 12 663
rect -12 458 -9 657
rect 9 458 12 657
rect -12 452 12 458
rect -12 -458 12 -452
rect -12 -657 -9 -458
rect 9 -657 12 -458
rect -12 -663 12 -657
<< res0p35 >>
rect -18 -451 18 451
<< properties >>
string FIXED_BBOX -74 -722 74 722
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 9.0 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 52.504k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
