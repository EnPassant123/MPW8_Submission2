magic
tech sky130A
magscale 1 2
timestamp 1672468335
<< metal3 >>
rect -5454 5134 -120 5162
rect -5454 148 -204 5134
rect -140 148 -120 5134
rect -5454 120 -120 148
rect 120 5134 5454 5162
rect 120 148 5370 5134
rect 5434 148 5454 5134
rect 120 120 5454 148
rect -5454 -148 -120 -120
rect -5454 -5134 -204 -148
rect -140 -5134 -120 -148
rect -5454 -5162 -120 -5134
rect 120 -148 5454 -120
rect 120 -5134 5370 -148
rect 5434 -5134 5454 -148
rect 120 -5162 5454 -5134
<< via3 >>
rect -204 148 -140 5134
rect 5370 148 5434 5134
rect -204 -5134 -140 -148
rect 5370 -5134 5434 -148
<< mimcap >>
rect -5414 5082 -452 5122
rect -5414 200 -5374 5082
rect -492 200 -452 5082
rect -5414 160 -452 200
rect 160 5082 5122 5122
rect 160 200 200 5082
rect 5082 200 5122 5082
rect 160 160 5122 200
rect -5414 -200 -452 -160
rect -5414 -5082 -5374 -200
rect -492 -5082 -452 -200
rect -5414 -5122 -452 -5082
rect 160 -200 5122 -160
rect 160 -5082 200 -200
rect 5082 -5082 5122 -200
rect 160 -5122 5122 -5082
<< mimcapcontact >>
rect -5374 200 -492 5082
rect 200 200 5082 5082
rect -5374 -5082 -492 -200
rect 200 -5082 5082 -200
<< metal4 >>
rect -2985 5083 -2881 5282
rect -224 5134 -120 5282
rect -5375 5082 -491 5083
rect -5375 200 -5374 5082
rect -492 200 -491 5082
rect -5375 199 -491 200
rect -2985 -199 -2881 199
rect -224 148 -204 5134
rect -140 148 -120 5134
rect 2589 5083 2693 5282
rect 5350 5134 5454 5282
rect 199 5082 5083 5083
rect 199 200 200 5082
rect 5082 200 5083 5082
rect 199 199 5083 200
rect -224 -148 -120 148
rect -5375 -200 -491 -199
rect -5375 -5082 -5374 -200
rect -492 -5082 -491 -200
rect -5375 -5083 -491 -5082
rect -2985 -5282 -2881 -5083
rect -224 -5134 -204 -148
rect -140 -5134 -120 -148
rect 2589 -199 2693 199
rect 5350 148 5370 5134
rect 5434 148 5454 5134
rect 5350 -148 5454 148
rect 199 -200 5083 -199
rect 199 -5082 200 -200
rect 5082 -5082 5083 -200
rect 199 -5083 5083 -5082
rect -224 -5282 -120 -5134
rect 2589 -5282 2693 -5083
rect 5350 -5134 5370 -148
rect 5434 -5134 5454 -148
rect 5350 -5282 5454 -5134
<< properties >>
string FIXED_BBOX 120 120 5162 5162
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 24.805 l 24.805 val 1.249k carea 2.00 cperi 0.19 nx 2 ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
