magic
tech sky130A
magscale 1 2
timestamp 1672354625
<< error_p >>
rect -29 1072 29 1078
rect -29 1038 -17 1072
rect -29 1032 29 1038
rect -29 -1038 29 -1032
rect -29 -1072 -17 -1038
rect -29 -1078 29 -1072
<< pwell >>
rect -212 -1210 212 1210
<< nmoslvt >>
rect -16 -1000 16 1000
<< ndiff >>
rect -74 988 -16 1000
rect -74 -988 -62 988
rect -28 -988 -16 988
rect -74 -1000 -16 -988
rect 16 988 74 1000
rect 16 -988 28 988
rect 62 -988 74 988
rect 16 -1000 74 -988
<< ndiffc >>
rect -62 -988 -28 988
rect 28 -988 62 988
<< psubdiff >>
rect -176 1140 -80 1174
rect 80 1140 176 1174
rect -176 1078 -142 1140
rect 142 1078 176 1140
rect -176 -1140 -142 -1078
rect 142 -1140 176 -1078
rect -176 -1174 -80 -1140
rect 80 -1174 176 -1140
<< psubdiffcont >>
rect -80 1140 80 1174
rect -176 -1078 -142 1078
rect 142 -1078 176 1078
rect -80 -1174 80 -1140
<< poly >>
rect -33 1072 33 1088
rect -33 1038 -17 1072
rect 17 1038 33 1072
rect -33 1022 33 1038
rect -16 1000 16 1022
rect -16 -1022 16 -1000
rect -33 -1038 33 -1022
rect -33 -1072 -17 -1038
rect 17 -1072 33 -1038
rect -33 -1088 33 -1072
<< polycont >>
rect -17 1038 17 1072
rect -17 -1072 17 -1038
<< locali >>
rect -176 1140 -80 1174
rect 80 1140 176 1174
rect -176 1078 -142 1140
rect 142 1078 176 1140
rect -33 1038 -17 1072
rect 17 1038 33 1072
rect -62 988 -28 1004
rect -62 -1004 -28 -988
rect 28 988 62 1004
rect 28 -1004 62 -988
rect -33 -1072 -17 -1038
rect 17 -1072 33 -1038
rect -176 -1140 -142 -1078
rect 142 -1140 176 -1078
rect -176 -1174 -80 -1140
rect 80 -1174 176 -1140
<< viali >>
rect -17 1038 17 1072
rect -62 -988 -28 988
rect 28 -988 62 988
rect -17 -1072 17 -1038
<< metal1 >>
rect -29 1072 29 1078
rect -29 1038 -17 1072
rect 17 1038 29 1072
rect -29 1032 29 1038
rect -68 988 -22 1000
rect -68 -988 -62 988
rect -28 -988 -22 988
rect -68 -1000 -22 -988
rect 22 988 68 1000
rect 22 -988 28 988
rect 62 -988 68 988
rect 22 -1000 68 -988
rect -29 -1038 29 -1032
rect -29 -1072 -17 -1038
rect 17 -1072 29 -1038
rect -29 -1078 29 -1072
<< properties >>
string FIXED_BBOX -159 -1157 159 1157
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 10.0 l 0.155 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
