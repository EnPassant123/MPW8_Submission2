magic
tech sky130A
magscale 1 2
timestamp 1672366060
<< locali >>
rect -3475 2439 -745 2445
rect -3475 2401 -2229 2439
rect -2191 2401 -745 2439
rect -3475 2365 -745 2401
rect -2105 1109 -1655 1115
rect -2105 1071 -1699 1109
rect -1661 1071 -1655 1109
rect -2105 1065 -1655 1071
rect -4085 935 -2255 985
rect -2305 705 -2255 935
rect -2105 885 -2055 1065
rect -1915 945 105 995
rect -1915 705 -1865 945
rect -2305 655 -1865 705
rect -125 -226 -75 -220
rect -125 -264 -119 -226
rect -81 -264 -75 -226
rect -125 -465 -75 -264
rect -4275 -515 -75 -465
rect 55 -615 105 945
rect -1185 -665 105 -615
rect -3255 -1605 -3205 -705
rect -1185 -1605 -1135 -665
rect -3255 -1655 -1135 -1605
rect -3255 -2875 -3205 -1655
rect -1875 -1796 -1825 -1655
rect -1875 -1834 -1869 -1796
rect -1831 -1834 -1825 -1796
rect -1875 -1840 -1825 -1834
rect -1185 -2895 -1135 -1655
<< viali >>
rect -2229 2401 -2191 2439
rect -1699 1071 -1661 1109
rect -2105 835 -2055 885
rect -119 -264 -81 -226
rect -4325 -515 -4275 -465
rect -1869 -1834 -1831 -1796
<< metal1 >>
rect -2235 2439 -2185 2451
rect -2235 2401 -2229 2439
rect -2191 2401 -2185 2439
rect -3400 2260 -3300 2310
rect -2235 2210 -2185 2401
rect -1000 2260 -900 2310
rect -1100 2210 -1000 2220
rect -3510 2160 -3410 2210
rect -3295 2170 -1000 2210
rect -3295 2160 -1015 2170
rect -900 2160 -800 2210
rect -3465 1455 -3415 2160
rect -3865 1405 -3415 1455
rect -3295 1425 -3245 2160
rect -1065 1435 -1015 2160
rect -895 1485 -845 2160
rect -895 1435 -585 1485
rect -3865 1175 -3815 1405
rect -3400 1330 -895 1380
rect -4285 1125 -1855 1175
rect -4285 810 -4235 1125
rect -4030 840 -3930 890
rect -2830 840 -2730 890
rect -2117 885 -2043 891
rect -2395 835 -2105 885
rect -2055 835 -2043 885
rect -4285 760 -4010 810
rect -3965 760 -3860 810
rect -2910 760 -2810 810
rect -2760 805 -2660 810
rect -2395 805 -2345 835
rect -2117 829 -2043 835
rect -3965 -135 -3915 760
rect -2865 -135 -2815 760
rect -3965 -185 -2815 -135
rect -2765 755 -2345 805
rect -1905 815 -1855 1125
rect -635 1115 -585 1435
rect -1711 1109 -115 1115
rect -1711 1071 -1699 1109
rect -1661 1071 -115 1109
rect -1711 1065 -115 1071
rect -1630 840 -1530 890
rect -440 840 -340 890
rect -1905 810 -1711 815
rect -165 810 -115 1065
rect -1905 765 -1610 810
rect -1801 760 -1610 765
rect -1565 760 -1460 810
rect -510 760 -410 810
rect -365 760 -115 810
rect -4050 -225 -3950 -220
rect -4325 -270 -3950 -225
rect -4325 -275 -3955 -270
rect -4325 -453 -4275 -275
rect -4331 -465 -4269 -453
rect -4331 -515 -4325 -465
rect -4275 -515 -4269 -465
rect -4331 -527 -4269 -515
rect -3615 -789 -3565 -185
rect -2765 -190 -2715 755
rect -1665 -190 -1615 760
rect -1565 -135 -1515 760
rect -465 -135 -415 760
rect -1565 -185 -415 -135
rect -365 -185 -315 760
rect -2850 -270 -1535 -220
rect -1640 -280 -1540 -270
rect -3430 -760 -3330 -710
rect -1050 -760 -950 -710
rect -3615 -795 -3419 -789
rect -3615 -845 -3415 -795
rect -1065 -800 -1015 -795
rect -775 -800 -725 -185
rect -440 -226 -69 -220
rect -440 -264 -119 -226
rect -81 -264 -69 -226
rect -440 -270 -69 -264
rect -3520 -850 -3419 -845
rect -3469 -2779 -3419 -850
rect -3365 -850 -3260 -800
rect -1110 -850 -1010 -800
rect -960 -850 -725 -800
rect -3365 -2733 -3309 -850
rect -2565 -1475 -1585 -1425
rect -2565 -1795 -2515 -1475
rect -2240 -1760 -2140 -1710
rect -2565 -1800 -2215 -1795
rect -2170 -1796 -1805 -1790
rect -2565 -1845 -2210 -1800
rect -2170 -1834 -1869 -1796
rect -1831 -1834 -1805 -1796
rect -2170 -1840 -1805 -1834
rect -2310 -1850 -2210 -1845
rect -3365 -2735 -2969 -2733
rect -2265 -2735 -2215 -1850
rect -3365 -2785 -2215 -2735
rect -2163 -2785 -2113 -1840
rect -1635 -2735 -1585 -1475
rect -1065 -2735 -1015 -850
rect -1635 -2785 -1015 -2735
rect -957 -2783 -907 -850
rect -3735 -2870 -3340 -2820
rect -2240 -2870 -1745 -2820
rect -1040 -2870 -705 -2820
use sky130_fd_pr__nfet_01v8_lvt_9DW9LC  XM7
timestamp 1672366060
transform 1 0 -3387 0 1 -1788
box -212 -1210 212 1210
use sky130_fd_pr__nfet_01v8_lvt_84HFGD  XM9
timestamp 1672366060
transform 1 0 -1587 0 1 312
box -212 -710 212 710
use sky130_fd_pr__nfet_01v8_lvt_84HFGD  XM10
timestamp 1672366060
transform 1 0 -387 0 1 312
box -212 -710 212 710
use sky130_fd_pr__nfet_01v8_lvt_84HFGD  XM11
timestamp 1672366060
transform 1 0 -2787 0 1 312
box -212 -710 212 710
use sky130_fd_pr__nfet_01v8_lvt_9DW9LC  sky130_fd_pr__nfet_01v8_lvt_9DW9LC_0
timestamp 1672366060
transform 1 0 -987 0 1 -1788
box -212 -1210 212 1210
use sky130_fd_pr__nfet_01v8_lvt_84HFGD  sky130_fd_pr__nfet_01v8_lvt_84HFGD_0
timestamp 1672366060
transform 1 0 -3987 0 1 312
box -212 -710 212 710
use sky130_fd_pr__nfet_01v8_lvt_84HFGD  sky130_fd_pr__nfet_01v8_lvt_84HFGD_1
timestamp 1672366060
transform 1 0 -2187 0 1 -2288
box -212 -710 212 710
use sky130_fd_pr__pfet_01v8_lvt_NK53LE  sky130_fd_pr__pfet_01v8_lvt_NK53LE_0
timestamp 1672366060
transform 1 0 -3352 0 1 1819
box -247 -619 247 619
use sky130_fd_pr__pfet_01v8_lvt_NK53LE  sky130_fd_pr__pfet_01v8_lvt_NK53LE_1
timestamp 1672366060
transform 1 0 -952 0 1 1819
box -247 -619 247 619
<< labels >>
rlabel locali -2155 2365 -2105 2415 1 vcc
port 0 n
rlabel metal1 -4325 -405 -4275 -355 1 LO+
port 1 n
rlabel metal1 -2295 -270 -2245 -220 1 LO-
port 2 n
rlabel metal1 -3735 -2870 -3685 -2820 1 RF+
port 3 n
rlabel metal1 -755 -2870 -705 -2820 1 RF-
port 4 n
rlabel metal1 -3825 1125 -3775 1175 1 IF+
port 5 n
rlabel metal1 -1005 1065 -955 1115 1 IF-
port 6 n
rlabel metal1 -1835 -2870 -1785 -2820 1 NB
port 7 n
rlabel metal1 -2185 1330 -2135 1380 1 PB
port 8 n
rlabel metal1 -1945 -1840 -1895 -1790 1 GND
port 9 n
<< end >>
