magic
tech sky130A
magscale 1 2
timestamp 1672474592
<< metal3 >>
rect -2687 2513 2687 2541
rect -2687 -2513 2603 2513
rect 2667 -2513 2687 2513
rect -2687 -2541 2687 -2513
<< via3 >>
rect 2603 -2513 2667 2513
<< mimcap >>
rect -2647 2461 2355 2501
rect -2647 -2461 -2607 2461
rect 2315 -2461 2355 2461
rect -2647 -2501 2355 -2461
<< mimcapcontact >>
rect -2607 -2461 2315 2461
<< metal4 >>
rect 2587 2513 2683 2529
rect -2608 2461 2316 2462
rect -2608 -2461 -2607 2461
rect 2315 -2461 2316 2461
rect -2608 -2462 2316 -2461
rect 2587 -2513 2603 2513
rect 2667 -2513 2683 2513
rect 2587 -2529 2683 -2513
<< properties >>
string FIXED_BBOX -2687 -2541 2395 2541
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 25.005 l 25.005 val 1.269k carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
