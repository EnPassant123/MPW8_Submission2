magic
tech sky130A
timestamp 1606063140
<< pwell >>
rect -481 -229 481 229
<< mvnmos >>
rect -367 -100 -287 100
rect -258 -100 -178 100
rect -149 -100 -69 100
rect -40 -100 40 100
rect 69 -100 149 100
rect 178 -100 258 100
rect 287 -100 367 100
<< mvndiff >>
rect -396 94 -367 100
rect -396 -94 -390 94
rect -373 -94 -367 94
rect -396 -100 -367 -94
rect -287 94 -258 100
rect -287 -94 -281 94
rect -264 -94 -258 94
rect -287 -100 -258 -94
rect -178 94 -149 100
rect -178 -94 -172 94
rect -155 -94 -149 94
rect -178 -100 -149 -94
rect -69 94 -40 100
rect -69 -94 -63 94
rect -46 -94 -40 94
rect -69 -100 -40 -94
rect 40 94 69 100
rect 40 -94 46 94
rect 63 -94 69 94
rect 40 -100 69 -94
rect 149 94 178 100
rect 149 -94 155 94
rect 172 -94 178 94
rect 149 -100 178 -94
rect 258 94 287 100
rect 258 -94 264 94
rect 281 -94 287 94
rect 258 -100 287 -94
rect 367 94 396 100
rect 367 -94 373 94
rect 390 -94 396 94
rect 367 -100 396 -94
<< mvndiffc >>
rect -390 -94 -373 94
rect -281 -94 -264 94
rect -172 -94 -155 94
rect -63 -94 -46 94
rect 46 -94 63 94
rect 155 -94 172 94
rect 264 -94 281 94
rect 373 -94 390 94
<< mvpsubdiff >>
rect -463 205 463 211
rect -463 188 -409 205
rect 409 188 463 205
rect -463 182 463 188
rect -463 157 -434 182
rect -463 -157 -457 157
rect -440 -157 -434 157
rect 434 157 463 182
rect -463 -182 -434 -157
rect 434 -157 440 157
rect 457 -157 463 157
rect 434 -182 463 -157
rect -463 -188 463 -182
rect -463 -205 -409 -188
rect 409 -205 463 -188
rect -463 -211 463 -205
<< mvpsubdiffcont >>
rect -409 188 409 205
rect -457 -157 -440 157
rect 440 -157 457 157
rect -409 -205 409 -188
<< poly >>
rect -367 136 -287 144
rect -367 119 -359 136
rect -295 119 -287 136
rect -367 100 -287 119
rect -258 136 -178 144
rect -258 119 -250 136
rect -186 119 -178 136
rect -258 100 -178 119
rect -149 136 -69 144
rect -149 119 -141 136
rect -77 119 -69 136
rect -149 100 -69 119
rect -40 136 40 144
rect -40 119 -32 136
rect 32 119 40 136
rect -40 100 40 119
rect 69 136 149 144
rect 69 119 77 136
rect 141 119 149 136
rect 69 100 149 119
rect 178 136 258 144
rect 178 119 186 136
rect 250 119 258 136
rect 178 100 258 119
rect 287 136 367 144
rect 287 119 295 136
rect 359 119 367 136
rect 287 100 367 119
rect -367 -119 -287 -100
rect -367 -136 -359 -119
rect -295 -136 -287 -119
rect -367 -144 -287 -136
rect -258 -119 -178 -100
rect -258 -136 -250 -119
rect -186 -136 -178 -119
rect -258 -144 -178 -136
rect -149 -119 -69 -100
rect -149 -136 -141 -119
rect -77 -136 -69 -119
rect -149 -144 -69 -136
rect -40 -119 40 -100
rect -40 -136 -32 -119
rect 32 -136 40 -119
rect -40 -144 40 -136
rect 69 -119 149 -100
rect 69 -136 77 -119
rect 141 -136 149 -119
rect 69 -144 149 -136
rect 178 -119 258 -100
rect 178 -136 186 -119
rect 250 -136 258 -119
rect 178 -144 258 -136
rect 287 -119 367 -100
rect 287 -136 295 -119
rect 359 -136 367 -119
rect 287 -144 367 -136
<< polycont >>
rect -359 119 -295 136
rect -250 119 -186 136
rect -141 119 -77 136
rect -32 119 32 136
rect 77 119 141 136
rect 186 119 250 136
rect 295 119 359 136
rect -359 -136 -295 -119
rect -250 -136 -186 -119
rect -141 -136 -77 -119
rect -32 -136 32 -119
rect 77 -136 141 -119
rect 186 -136 250 -119
rect 295 -136 359 -119
<< locali >>
rect -457 188 -409 205
rect 409 188 457 205
rect -457 157 -440 188
rect 440 157 457 188
rect -367 119 -359 136
rect -295 119 -287 136
rect -258 119 -250 136
rect -186 119 -178 136
rect -149 119 -141 136
rect -77 119 -69 136
rect -40 119 -32 136
rect 32 119 40 136
rect 69 119 77 136
rect 141 119 149 136
rect 178 119 186 136
rect 250 119 258 136
rect 287 119 295 136
rect 359 119 367 136
rect -390 94 -373 102
rect -390 -102 -373 -94
rect -281 94 -264 102
rect -281 -102 -264 -94
rect -172 94 -155 102
rect -172 -102 -155 -94
rect -63 94 -46 102
rect -63 -102 -46 -94
rect 46 94 63 102
rect 46 -102 63 -94
rect 155 94 172 102
rect 155 -102 172 -94
rect 264 94 281 102
rect 264 -102 281 -94
rect 373 94 390 102
rect 373 -102 390 -94
rect -367 -136 -359 -119
rect -295 -136 -287 -119
rect -258 -136 -250 -119
rect -186 -136 -178 -119
rect -149 -136 -141 -119
rect -77 -136 -69 -119
rect -40 -136 -32 -119
rect 32 -136 40 -119
rect 69 -136 77 -119
rect 141 -136 149 -119
rect 178 -136 186 -119
rect 250 -136 258 -119
rect 287 -136 295 -119
rect 359 -136 367 -119
rect -457 -188 -440 -157
rect 440 -188 457 -157
rect -457 -205 -409 -188
rect 409 -205 457 -188
<< viali >>
rect -457 -131 -440 131
rect -359 119 -295 136
rect -250 119 -186 136
rect -141 119 -77 136
rect -32 119 32 136
rect 77 119 141 136
rect 186 119 250 136
rect 295 119 359 136
rect -390 10 -373 85
rect -281 -85 -264 -10
rect -172 10 -155 85
rect -63 -85 -46 -10
rect 46 10 63 85
rect 155 -85 172 -10
rect 264 10 281 85
rect 373 -85 390 -10
rect -359 -136 -295 -119
rect -250 -136 -186 -119
rect -141 -136 -77 -119
rect -32 -136 32 -119
rect 77 -136 141 -119
rect 186 -136 250 -119
rect 295 -136 359 -119
<< metal1 >>
rect -460 131 -437 137
rect -460 -131 -457 131
rect -440 -131 -437 131
rect -365 136 -289 139
rect -365 119 -359 136
rect -295 119 -289 136
rect -365 116 -289 119
rect -256 136 -180 139
rect -256 119 -250 136
rect -186 119 -180 136
rect -256 116 -180 119
rect -147 136 -71 139
rect -147 119 -141 136
rect -77 119 -71 136
rect -147 116 -71 119
rect -38 136 38 139
rect -38 119 -32 136
rect 32 119 38 136
rect -38 116 38 119
rect 71 136 147 139
rect 71 119 77 136
rect 141 119 147 136
rect 71 116 147 119
rect 180 136 256 139
rect 180 119 186 136
rect 250 119 256 136
rect 180 116 256 119
rect 289 136 365 139
rect 289 119 295 136
rect 359 119 365 136
rect 289 116 365 119
rect -393 85 -370 91
rect -393 10 -390 85
rect -373 10 -370 85
rect -393 4 -370 10
rect -175 85 -152 91
rect -175 10 -172 85
rect -155 10 -152 85
rect -175 4 -152 10
rect 43 85 66 91
rect 43 10 46 85
rect 63 10 66 85
rect 43 4 66 10
rect 261 85 284 91
rect 261 10 264 85
rect 281 10 284 85
rect 261 4 284 10
rect -284 -10 -261 -4
rect -284 -85 -281 -10
rect -264 -85 -261 -10
rect -284 -91 -261 -85
rect -66 -10 -43 -4
rect -66 -85 -63 -10
rect -46 -85 -43 -10
rect -66 -91 -43 -85
rect 152 -10 175 -4
rect 152 -85 155 -10
rect 172 -85 175 -10
rect 152 -91 175 -85
rect 370 -10 393 -4
rect 370 -85 373 -10
rect 390 -85 393 -10
rect 370 -91 393 -85
rect -460 -137 -437 -131
rect -365 -119 -289 -116
rect -365 -136 -359 -119
rect -295 -136 -289 -119
rect -365 -139 -289 -136
rect -256 -119 -180 -116
rect -256 -136 -250 -119
rect -186 -136 -180 -119
rect -256 -139 -180 -136
rect -147 -119 -71 -116
rect -147 -136 -141 -119
rect -77 -136 -71 -119
rect -147 -139 -71 -136
rect -38 -119 38 -116
rect -38 -136 -32 -119
rect 32 -136 38 -119
rect -38 -139 38 -136
rect 71 -119 147 -116
rect 71 -136 77 -119
rect 141 -136 147 -119
rect 71 -139 147 -136
rect 180 -119 256 -116
rect 180 -136 186 -119
rect 250 -136 256 -119
rect 180 -139 256 -136
rect 289 -119 365 -116
rect 289 -136 295 -119
rect 359 -136 365 -119
rect 289 -139 365 -136
<< properties >>
string FIXED_BBOX -448 -196 448 196
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 2.00 l 0.80 m 1 nf 7 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc +40 viadrn -40 viagate 100 viagb 0 viagr 0 viagl 70 viagt 0
<< end >>
