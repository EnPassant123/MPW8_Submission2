magic
tech sky130A
timestamp 1671954411
<< metal3 >>
rect -1343 1256 1343 1270
rect -1343 -1256 1301 1256
rect 1333 -1256 1343 1256
rect -1343 -1270 1343 -1256
<< via3 >>
rect 1301 -1256 1333 1256
<< mimcap >>
rect -1323 1230 1177 1250
rect -1323 -1230 -1303 1230
rect 1157 -1230 1177 1230
rect -1323 -1250 1177 -1230
<< mimcapcontact >>
rect -1303 -1230 1157 1230
<< metal4 >>
rect 1293 1256 1341 1264
rect 1293 -1256 1301 1256
rect 1333 -1256 1341 1256
rect 1293 -1264 1341 -1256
<< properties >>
string FIXED_BBOX -1343 -1270 1197 1270
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 25 l 25 val 1.269k carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
