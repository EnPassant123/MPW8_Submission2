magic
tech sky130A
timestamp 1671945152
<< metal3 >>
rect -843 756 843 770
rect -843 -756 801 756
rect 833 -756 843 756
rect -843 -770 843 -756
<< via3 >>
rect 801 -756 833 756
<< mimcap >>
rect -823 730 677 750
rect -823 -730 -803 730
rect 657 -730 677 730
rect -823 -750 677 -730
<< mimcapcontact >>
rect -803 -730 657 730
<< metal4 >>
rect 793 756 841 764
rect 793 -756 801 756
rect 833 -756 841 756
rect 793 -764 841 -756
<< properties >>
string FIXED_BBOX -843 -770 697 770
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 15 l 15 val 461.4 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
