magic
tech sky130A
magscale 1 2
timestamp 1672362834
<< metal3 >>
rect -3186 3012 3186 3040
rect -3186 -3012 3102 3012
rect 3166 -3012 3186 3012
rect -3186 -3040 3186 -3012
<< via3 >>
rect 3102 -3012 3166 3012
<< mimcap >>
rect -3146 2960 2854 3000
rect -3146 -2960 -3106 2960
rect 2814 -2960 2854 2960
rect -3146 -3000 2854 -2960
<< mimcapcontact >>
rect -3106 -2960 2814 2960
<< metal4 >>
rect 3086 3012 3182 3028
rect -3107 2960 2815 2961
rect -3107 -2960 -3106 2960
rect 2814 -2960 2815 2960
rect -3107 -2961 2815 -2960
rect 3086 -3012 3102 3012
rect 3166 -3012 3182 3012
rect 3086 -3028 3182 -3012
<< properties >>
string FIXED_BBOX -3186 -3040 2894 3040
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 29.995 l 29.995 val 1.822k carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
