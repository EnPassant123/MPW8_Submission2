magic
tech sky130A
magscale 1 2
timestamp 1672466235
<< metal3 >>
rect -1587 1413 1587 1441
rect -1587 -1413 1503 1413
rect 1567 -1413 1587 1413
rect -1587 -1441 1587 -1413
<< via3 >>
rect 1503 -1413 1567 1413
<< mimcap >>
rect -1547 1361 1255 1401
rect -1547 -1361 -1507 1361
rect 1215 -1361 1255 1361
rect -1547 -1401 1255 -1361
<< mimcapcontact >>
rect -1507 -1361 1215 1361
<< metal4 >>
rect 1487 1413 1583 1429
rect -1508 1361 1216 1362
rect -1508 -1361 -1507 1361
rect 1215 -1361 1216 1361
rect -1508 -1362 1216 -1361
rect 1487 -1413 1503 1413
rect 1567 -1413 1583 1413
rect 1487 -1429 1583 -1413
<< properties >>
string FIXED_BBOX -1587 -1441 1295 1441
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 14.005 l 14.005 val 402.923 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
