* NGSPICE file created from user_analog_project_wrapper.ext - technology: sky130A

.subckt sky130_fd_pr__cap_mim_m3_1_P68BUM m3_n3186_n3040# c1_n3146_n3000#
X0 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_PH9SS5 a_n50_n297# a_50_n200# a_n108_n200# w_n246_n419#
X0 a_50_n200# a_n50_n297# a_n108_n200# w_n246_n419# sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_SMGWK2 a_n210_n574# a_50_n400# a_n108_n400# a_n50_n488#
X0 a_50_n400# a_n50_n488# a_n108_n400# a_n210_n574# sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
.ends

.subckt analogsub vdd Vplus voffset Vminus Nbias vout gnd
Xsky130_fd_pr__pfet_01v8_lvt_PH9SS5_0 m1_n1210_2130# m1_n1210_2130# vdd vdd sky130_fd_pr__pfet_01v8_lvt_PH9SS5
Xsky130_fd_pr__pfet_01v8_lvt_PH9SS5_1 m1_n1210_2130# vdd vout vdd sky130_fd_pr__pfet_01v8_lvt_PH9SS5
Xsky130_fd_pr__pfet_01v8_lvt_PH9SS5_2 m1_391_2121# vout vdd vdd sky130_fd_pr__pfet_01v8_lvt_PH9SS5
Xsky130_fd_pr__pfet_01v8_lvt_PH9SS5_3 m1_391_2121# vdd m1_391_2121# vdd sky130_fd_pr__pfet_01v8_lvt_PH9SS5
XXM112 gnd vout m1_0_490# Vminus sky130_fd_pr__nfet_01v8_lvt_SMGWK2
XXM113 gnd m1_0_490# m1_391_2121# Vplus sky130_fd_pr__nfet_01v8_lvt_SMGWK2
XXM114 gnd gnd m1_0_490# Nbias sky130_fd_pr__nfet_01v8_lvt_SMGWK2
XXM117 gnd m1_n1210_2130# m1_n1330_400# voffset sky130_fd_pr__nfet_01v8_lvt_SMGWK2
XXM118 gnd m1_n1330_400# vout vout sky130_fd_pr__nfet_01v8_lvt_SMGWK2
XXM119 gnd gnd m1_n1330_400# Nbias sky130_fd_pr__nfet_01v8_lvt_SMGWK2
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_R9FY7S a_n35_n1483# a_n35_1051# a_n165_n1613#
X0 a_n35_n1483# a_n35_1051# a_n165_n1613# sky130_fd_pr__res_xhigh_po_0p35 l=1.051e+07u
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_REKGFF m3_n2687_n2541# c1_n2647_n2501#
X0 c1_n2647_n2501# m3_n2687_n2541# sky130_fd_pr__cap_mim_m3_1 l=2.501e+07u w=2.501e+07u
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_5B6GLN c1_n1647_n1501# m3_n1687_n1541#
X0 c1_n1647_n1501# m3_n1687_n1541# sky130_fd_pr__cap_mim_m3_1 l=1.501e+07u w=1.501e+07u
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VPWR X VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=9.1e+11p pd=7.82e+06u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=3.801e+11p pd=4.33e+06u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfrbp_1 CLK D RESET_B VGND VPWR Q Q_N VNB VPB
X0 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=1.5393e+12p ps=1.452e+07u w=1e+06u l=150000u
X1 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X2 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X3 VPWR a_1283_21# a_1847_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X4 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X5 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X6 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X7 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=1.2225e+12p pd=1.139e+07u as=0p ps=0u w=420000u l=150000u
X8 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X9 Q_N a_1847_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X10 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X11 VGND a_1283_21# a_1847_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X12 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X16 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X17 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X21 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X22 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X24 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X27 Q_N a_1847_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X28 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X31 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_1 A VGND VPWR Y VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.268e+11p pd=2.22e+06u as=4.536e+11p ps=4.44e+06u w=840000u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=1.197e+11p pd=1.41e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt quadgen clkin outa outb outc outd sky130_fd_sc_hd__tapvpwrvgnd_1_2/VPWR gnd
+ vcc sky130_fd_sc_hd__tapvpwrvgnd_1_2/VGND
Xsky130_fd_sc_hd__clkbuf_4_0 x10/Q_N gnd vcc outc gnd vcc sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_1 x10/Q gnd vcc outd gnd vcc sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_2 sky130_fd_sc_hd__clkbuf_4_2/A gnd vcc outb gnd vcc sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_4_3 x10/D gnd vcc outa gnd vcc sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__dfrbp_1_0 clkin x10/Q_N vcc gnd vcc x10/D sky130_fd_sc_hd__clkbuf_4_2/A
+ gnd vcc sky130_fd_sc_hd__dfrbp_1
Xx10 x33/Y x10/D vcc gnd vcc x10/Q x10/Q_N gnd vcc sky130_fd_sc_hd__dfrbp_1
Xx33 clkin gnd vcc x33/Y gnd vcc sky130_fd_sc_hd__clkinv_1
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_U9BGXT a_n108_n300# a_n50_n388# a_n210_n474# a_50_n300#
X0 a_50_n300# a_n50_n388# a_n108_n300# a_n210_n474# sky130_fd_pr__nfet_01v8_lvt ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=500000u
.ends

.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VPWR X VNB VPB
X0 VGND A a_311_413# VNB sky130_fd_pr__nfet_01v8 ad=5.5025e+11p pd=6.15e+06u as=2.331e+11p ps=2.79e+06u w=420000u l=150000u
X1 VPWR A a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=5.41725e+11p pd=5.32e+06u as=1.197e+11p ps=1.41e+06u w=420000u l=150000u
X2 a_393_413# a_205_93# a_311_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.43e+11p pd=2.66e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3 VGND C_N a_27_410# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4 VPWR C_N a_27_410# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5 X a_311_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.75e+11p pd=2.55e+06u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_27_410# a_311_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_561_297# B a_489_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X8 a_205_93# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X9 a_205_93# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X10 a_489_297# a_27_410# a_393_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_311_413# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_311_413# a_205_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 X a_311_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
.ends

.subckt clkdiv input output sky130_fd_sc_hd__tapvpwrvgnd_1_4/VPWR sky130_fd_sc_hd__tapvpwrvgnd_1_1/VPWR
+ x6/D x7/D sky130_fd_sc_hd__tapvpwrvgnd_1_2/VPWR vcc x5/D gnd
Xx5 input x5/D x7/RESET_B gnd vcc x5/Q x5/D gnd vcc sky130_fd_sc_hd__dfrbp_1
Xx6 x5/Q x6/D x7/RESET_B gnd vcc x6/Q x6/D gnd vcc sky130_fd_sc_hd__dfrbp_1
Xx7 x6/Q x7/D x7/RESET_B gnd vcc x7/Q x7/D gnd vcc sky130_fd_sc_hd__dfrbp_1
Xsky130_fd_sc_hd__or4bb_1_0 x5/D x6/D output x7/D gnd vcc x7/RESET_B gnd vcc sky130_fd_sc_hd__or4bb_1
Xsky130_fd_sc_hd__dfrbp_1_0 x7/Q output x7/RESET_B gnd vcc sky130_fd_sc_hd__dfrbp_1_0/Q
+ output gnd vcc sky130_fd_sc_hd__dfrbp_1
.ends

.subckt sky130_fd_pr__res_xhigh_po_5p73_WAQYE6 a_n573_516# a_n703_n1078# a_n573_n948#
X0 a_n573_n948# a_n573_516# a_n703_n1078# sky130_fd_pr__res_xhigh_po_5p73 l=5.16e+06u
.ends

.subckt sky130_fd_sc_hd__bufbuf_8 A VGND VPWR X VNB VPB
X0 a_318_47# a_206_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=5.3e+11p pd=5.06e+06u as=1.918e+12p ps=1.789e+07u w=1e+06u l=150000u
X1 VPWR a_318_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X2 VPWR a_206_47# a_318_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_318_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=7.02e+11p pd=7.36e+06u as=1.247e+12p ps=1.299e+07u w=650000u l=150000u
X4 X a_318_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR a_318_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X a_318_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND a_206_47# a_318_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X8 VPWR a_318_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_318_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_318_47# a_206_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X a_318_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_206_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X13 X a_318_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_206_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR a_318_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND a_206_47# a_318_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND a_318_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND a_318_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 VGND a_318_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 X a_318_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VGND a_318_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 VPWR a_206_47# a_318_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X24 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X25 X a_318_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkdlybuf4s50_1 A VGND VPWR X VNB VPB
X0 a_283_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=6.517e+11p ps=5.37e+06u w=820000u l=500000u
X1 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2 VPWR a_283_47# a_390_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X3 VGND a_283_47# a_390_47# VNB sky130_fd_pr__nfet_01v8 ad=4.027e+11p pd=3.97e+06u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X4 X a_390_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X6 a_283_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X7 X a_390_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_QP79FH a_n74_n1000# w_n212_n1219# a_n33_n1097# a_16_n1000#
X0 a_16_n1000# a_n33_n1097# a_n74_n1000# w_n212_n1219# sky130_fd_pr__pfet_01v8 ad=2.9e+12p pd=2.058e+07u as=2.9e+12p ps=2.058e+07u w=1e+07u l=160000u
.ends

.subckt sky130_fd_pr__nfet_01v8_A5ES5P a_n73_n1000# a_15_n1000# a_n33_n1088# a_n175_n1174#
X0 a_15_n1000# a_n33_n1088# a_n73_n1000# a_n175_n1174# sky130_fd_pr__nfet_01v8 ad=2.9e+12p pd=2.058e+07u as=2.9e+12p ps=2.058e+07u w=1e+07u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2_1 A B VGND VPWR Y VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=5.2e+11p pd=5.04e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt phasecmp a b out sky130_fd_sc_hd__tapvpwrvgnd_1_1/VPWR sky130_fd_sc_hd__tapvpwrvgnd_1_2/VGND
+ VSUBS vcc
XXR17 out VSUBS m1_5220_n910# sky130_fd_pr__res_xhigh_po_5p73_WAQYE6
Xx30 x39/B VSUBS vcc x30/X VSUBS vcc sky130_fd_sc_hd__bufbuf_8
Xx31 x39/Y VSUBS vcc x31/X VSUBS vcc sky130_fd_sc_hd__clkdlybuf4s50_1
XXM108 m1_5220_n910# vcc x162/X vcc sky130_fd_pr__pfet_01v8_QP79FH
XXM109 m1_5220_n910# VSUBS x30/X VSUBS sky130_fd_pr__nfet_01v8_A5ES5P
Xx28 b x31/X x31/X VSUBS vcc x39/B x28/Q_N VSUBS vcc sky130_fd_sc_hd__dfrbp_1
Xx39 x39/A x39/B VSUBS vcc x39/Y VSUBS vcc sky130_fd_sc_hd__nand2_1
Xx29 a x31/X x31/X VSUBS vcc x39/A x162/A VSUBS vcc sky130_fd_sc_hd__dfrbp_1
Xx162 x162/A VSUBS vcc x162/X VSUBS vcc sky130_fd_sc_hd__bufbuf_8
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_LU79P3 a_n35_n1303# a_n35_871# a_n165_n1433#
X0 a_n35_n1303# a_n35_871# a_n165_n1433# sky130_fd_pr__res_xhigh_po_0p35 l=8.71e+06u
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_PUMBUM m3_n6492_n12520# c1_n6452_n12480# c1_n13064_n12480#
+ m3_6732_n12520# c1_160_n12480# m3_120_n12520# m3_n13104_n12520# c1_6772_n12480#
X0 c1_n6452_n12480# m3_n6492_n12520# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X1 c1_n13064_n12480# m3_n13104_n12520# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X2 c1_6772_n12480# m3_6732_n12520# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X3 c1_n13064_n12480# m3_n13104_n12520# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X4 c1_n6452_n12480# m3_n6492_n12520# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X5 c1_6772_n12480# m3_6732_n12520# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X6 c1_n13064_n12480# m3_n13104_n12520# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X7 c1_160_n12480# m3_120_n12520# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X8 c1_6772_n12480# m3_6732_n12520# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X9 c1_160_n12480# m3_120_n12520# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X10 c1_160_n12480# m3_120_n12520# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X11 c1_n6452_n12480# m3_n6492_n12520# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X12 c1_n13064_n12480# m3_n13104_n12520# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X13 c1_160_n12480# m3_120_n12520# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X14 c1_6772_n12480# m3_6732_n12520# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X15 c1_n6452_n12480# m3_n6492_n12520# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_JDBWNB a_n108_n1000# a_50_n1000# a_n210_n1174#
+ a_n50_n1088#
X0 a_50_n1000# a_n50_n1088# a_n108_n1000# a_n210_n1174# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+12p pd=2.058e+07u as=2.9e+12p ps=2.058e+07u w=1e+07u l=500000u
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_R8KP6D c1_n5414_n5122# c1_160_n5122# m3_n5454_n5162#
+ m3_120_n5162#
X0 c1_160_n5122# m3_120_n5162# sky130_fd_pr__cap_mim_m3_1 l=2.481e+07u w=2.481e+07u
X1 c1_n5414_n5122# m3_n5454_n5162# sky130_fd_pr__cap_mim_m3_1 l=2.481e+07u w=2.481e+07u
X2 c1_n5414_n5122# m3_n5454_n5162# sky130_fd_pr__cap_mim_m3_1 l=2.481e+07u w=2.481e+07u
X3 c1_160_n5122# m3_120_n5162# sky130_fd_pr__cap_mim_m3_1 l=2.481e+07u w=2.481e+07u
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_G3F5X4 a_n35_3000# a_n165_n3562# a_n35_n3432#
X0 a_n35_n3432# a_n35_3000# a_n165_n3562# sky130_fd_pr__res_xhigh_po_0p35 l=3e+07u
.ends

.subckt sky130_fd_pr__res_xhigh_po_5p73_P7BAXV a_n573_n1433# a_n703_n1563# a_n573_1001#
X0 a_n573_n1433# a_n573_1001# a_n703_n1563# sky130_fd_pr__res_xhigh_po_5p73 l=1.001e+07u
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_TDASS5 a_n50_n597# a_50_n500# a_n108_n500# w_n246_n719#
X0 a_50_n500# a_n50_n597# a_n108_n500# w_n246_n719# sky130_fd_pr__pfet_01v8_lvt ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_X3MKZ5 a_n108_n1000# w_n246_n1219# a_n50_n1097#
+ a_50_n1000#
X0 a_50_n1000# a_n50_n1097# a_n108_n1000# w_n246_n1219# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+12p pd=2.058e+07u as=2.9e+12p ps=2.058e+07u w=1e+07u l=500000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_MYKW3H a_n50_n5988# a_n108_n5900# a_n210_n6074#
+ a_50_n5900#
X0 a_50_n5900# a_n50_n5988# a_n108_n5900# a_n210_n6074# sky130_fd_pr__nfet_01v8_lvt ad=1.711e+13p pd=1.1858e+08u as=1.711e+13p ps=1.1858e+08u w=5.9e+07u l=500000u
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_XP5BXZ a_n109_n300# w_n247_n519# a_n51_n397# a_51_n300#
X0 a_51_n300# a_n51_n397# a_n109_n300# w_n247_n519# sky130_fd_pr__pfet_01v8_lvt ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=510000u
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p69_FR2N8V a_n68_1040# a_n198_n1602# a_n68_n1472#
X0 a_n68_n1472# a_n68_1040# a_n198_n1602# sky130_fd_pr__res_xhigh_po_0p69 l=1.04e+07u
.ends

.subckt sky130_fd_pr__res_high_po_2p85_HV4VUF a_n284_1000# a_n284_n1432# a_n414_n1562#
X0 a_n284_n1432# a_n284_1000# a_n414_n1562# sky130_fd_pr__res_high_po_2p85 l=1e+07u
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_KYM84V m3_n886_n740# c1_n846_n700#
X0 c1_n846_n700# m3_n886_n740# sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_8TEW3F a_50_n500# a_n108_n500# a_n50_n588# a_n210_n674#
X0 a_50_n500# a_n50_n588# a_n108_n500# a_n210_n674# sky130_fd_pr__nfet_01v8_lvt ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_X3MVBA a_n108_n5000# w_n246_n5219# a_n50_n5097#
+ a_50_n5000#
X0 a_50_n5000# a_n50_n5097# a_n108_n5000# w_n246_n5219# sky130_fd_pr__pfet_01v8_lvt ad=1.45e+13p pd=1.0058e+08u as=1.45e+13p ps=1.0058e+08u w=5e+07u l=500000u
.ends

.subckt opamp vcc inv noninv output gnd
XXM56 m1_n2590_4110# vcc m1_n540_4980# vcc sky130_fd_pr__pfet_01v8_lvt_X3MKZ5
XXM57 li_1325_1915# output gnd gnd sky130_fd_pr__nfet_01v8_lvt_MYKW3H
XXM59 m1_n2580_3900# vcc m1_n540_3980# m1_n2590_4110# sky130_fd_pr__pfet_01v8_lvt_X3MKZ5
Xsky130_fd_pr__pfet_01v8_lvt_XP5BXZ_0 m1_n540_3980# vcc m1_n540_3980# m1_n540_4980#
+ sky130_fd_pr__pfet_01v8_lvt_XP5BXZ
Xsky130_fd_pr__pfet_01v8_lvt_XP5BXZ_1 m1_n2580_3900# vcc noninv li_1325_1915# sky130_fd_pr__pfet_01v8_lvt_XP5BXZ
XXR17 m1_n540_3980# gnd gnd sky130_fd_pr__res_xhigh_po_0p69_FR2N8V
XXR18 li_1325_1915# m1_3740_2320# gnd sky130_fd_pr__res_high_po_2p85_HV4VUF
XXC6 m1_3740_2320# output sky130_fd_pr__cap_mim_m3_1_KYM84V
XXM60 gnd m1_n2710_330# m1_n2710_330# gnd sky130_fd_pr__nfet_01v8_lvt_8TEW3F
XXM61 li_1325_1915# gnd m1_n2710_330# gnd sky130_fd_pr__nfet_01v8_lvt_8TEW3F
XXM62 vcc vcc m1_n540_4980# m1_1210_4110# sky130_fd_pr__pfet_01v8_lvt_X3MVBA
XXM63 m1_1210_4110# vcc m1_n540_3980# output sky130_fd_pr__pfet_01v8_lvt_X3MVBA
XXM53 m1_n540_4980# vcc m1_n540_4980# vcc sky130_fd_pr__pfet_01v8_lvt_XP5BXZ
XXM54 m1_n2710_330# vcc inv m1_n2580_3900# sky130_fd_pr__pfet_01v8_lvt_XP5BXZ
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_TE3E2R c1_n1547_n1401# m3_n1587_n1441#
X0 c1_n1547_n1401# m3_n1587_n1441# sky130_fd_pr__cap_mim_m3_1 l=1.401e+07u w=1.401e+07u
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p69_LVNRZ4 a_n68_690# a_n198_n1252# a_n68_n1122#
X0 a_n68_n1122# a_n68_690# a_n198_n1252# sky130_fd_pr__res_xhigh_po_0p69 l=6.9e+06u
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_4XRDQ9 a_n165_n1462# a_n35_900# a_n35_n1332#
X0 a_n35_n1332# a_n35_900# a_n165_n1462# sky130_fd_pr__res_xhigh_po_0p35 l=9e+06u
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_8R53B2 w_n247_n1219# a_n51_n1097# a_51_n1000#
+ a_n109_n1000#
X0 a_51_n1000# a_n51_n1097# a_n109_n1000# w_n247_n1219# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+12p pd=2.058e+07u as=2.9e+12p ps=2.058e+07u w=1e+07u l=510000u
.ends

.subckt sky130_fd_pr__res_xhigh_po_2p85_QPY2BD a_n284_950# a_n284_n1382# a_n414_n1512#
X0 a_n284_n1382# a_n284_950# a_n414_n1512# sky130_fd_pr__res_xhigh_po_2p85 l=9.5e+06u
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_NUYDZ7 c1_n3046_n9020# m3_n3086_n9060#
X0 c1_n3046_n9020# m3_n3086_n9060# sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=2.9e+07u
X1 c1_n3046_n9020# m3_n3086_n9060# sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=2.9e+07u
X2 c1_n3046_n9020# m3_n3086_n9060# sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=2.9e+07u
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_4BCNTW c1_n2146_n6160# m3_n2186_n6200#
X0 c1_n2146_n6160# m3_n2186_n6200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=2e+07u
X1 c1_n2146_n6160# m3_n2186_n6200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=2e+07u
.ends

.subckt filter vcc input out pb gnd
Xsky130_fd_pr__cap_mim_m3_1_TE3E2R_0 m1_19330_n37886# gnd sky130_fd_pr__cap_mim_m3_1_TE3E2R
XXR23 m1_20970_n34050# gnd m1_19330_n37886# sky130_fd_pr__res_xhigh_po_0p69_LVNRZ4
Xsky130_fd_pr__res_xhigh_po_0p35_4XRDQ9_0 gnd m1_21449_n33397# m1_20970_n34050# sky130_fd_pr__res_xhigh_po_0p35_4XRDQ9
Xsky130_fd_pr__pfet_01v8_lvt_8R53B2_0 vcc pb out vcc sky130_fd_pr__pfet_01v8_lvt_8R53B2
XXR7 m1_21449_n33397# input gnd sky130_fd_pr__res_xhigh_po_2p85_QPY2BD
XXC27 m1_21449_n33397# gnd sky130_fd_pr__cap_mim_m3_1_NUYDZ7
XXC4 out m1_20970_n34050# sky130_fd_pr__cap_mim_m3_1_4BCNTW
Xsky130_fd_pr__pfet_01v8_lvt_X3MKZ5_0 vcc m1_19330_n37886# gnd out sky130_fd_pr__pfet_01v8_lvt_8R53B2
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VPWR X VNB VPB
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.045e+12p pd=2.809e+07u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.24e+12p ps=2.048e+07u w=1e+06u l=150000u
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=1.2789e+12p ps=1.533e+07u w=420000u l=150000u
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.408e+11p ps=1.12e+07u w=420000u l=150000u
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_9DW9LC a_n74_n1000# a_16_n1000# a_n176_n1174#
+ a_n33_n1088#
X0 a_16_n1000# a_n33_n1088# a_n74_n1000# a_n176_n1174# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+12p pd=2.058e+07u as=2.9e+12p ps=2.058e+07u w=1e+07u l=160000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_84HFGD a_16_n500# a_n176_n674# a_n74_n500# a_n33_n588#
X0 a_16_n500# a_n33_n588# a_n74_n500# a_n176_n674# sky130_fd_pr__nfet_01v8_lvt ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=160000u
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_NK53LE w_n247_n619# a_n51_n497# a_51_n400# a_n109_n400#
X0 a_51_n400# a_n51_n497# a_n109_n400# w_n247_n619# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=510000u
.ends

.subckt gilbert vcc LO+ LO- RF+ RF- IF+ IF- NB PB GND
XXM7 m1_n3965_n185# m1_n3365_n2785# GND RF+ sky130_fd_pr__nfet_01v8_lvt_9DW9LC
XXM9 m1_n1565_n185# GND IF+ LO- sky130_fd_pr__nfet_01v8_lvt_84HFGD
Xsky130_fd_pr__pfet_01v8_lvt_NK53LE_0 vcc PB vcc IF+ sky130_fd_pr__pfet_01v8_lvt_NK53LE
Xsky130_fd_pr__nfet_01v8_lvt_84HFGD_0 m1_n3965_n185# GND IF+ LO+ sky130_fd_pr__nfet_01v8_lvt_84HFGD
Xsky130_fd_pr__pfet_01v8_lvt_NK53LE_1 vcc PB IF- vcc sky130_fd_pr__pfet_01v8_lvt_NK53LE
Xsky130_fd_pr__nfet_01v8_lvt_84HFGD_1 GND GND m1_n3365_n2785# NB sky130_fd_pr__nfet_01v8_lvt_84HFGD
Xsky130_fd_pr__nfet_01v8_lvt_9DW9LC_0 m1_n3365_n2785# m1_n1565_n185# GND RF- sky130_fd_pr__nfet_01v8_lvt_9DW9LC
XXM10 IF- GND m1_n1565_n185# LO+ sky130_fd_pr__nfet_01v8_lvt_84HFGD
XXM11 IF- GND m1_n3965_n185# LO- sky130_fd_pr__nfet_01v8_lvt_84HFGD
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_TRXTS5 a_n50_n597# a_50_n500# a_n108_n500# w_n246_n719#
X0 a_50_n500# a_n50_n597# a_n108_n500# w_n246_n719# sky130_fd_pr__pfet_01v8_lvt ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
.ends

.subckt sky130_fd_pr__nfet_01v8_Q8AFGD a_n74_n100# a_n33_n188# a_16_n100# a_n176_n274#
X0 a_16_n100# a_n33_n188# a_n74_n100# a_n176_n274# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=160000u
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_9SN4GA m3_n610_n464# c1_n570_n424#
X0 c1_n570_n424# m3_n610_n464# sky130_fd_pr__cap_mim_m3_1 l=4.24e+06u w=4.24e+06u
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VPWR X VNB VPB
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=2.291e+11p pd=2.16e+06u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=1.508e+11p ps=1.62e+06u w=520000u l=150000u
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_H4KU7R a_n35_1401# a_n165_n1963# a_n35_n1833#
X0 a_n35_n1833# a_n35_1401# a_n165_n1963# sky130_fd_pr__res_xhigh_po_0p35 l=1.401e+07u
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p69_ET3NLF a_n69_1231# a_n69_n1663# a_n199_n1793#
X0 a_n69_n1663# a_n69_1231# a_n199_n1793# sky130_fd_pr__res_xhigh_po_0p69 l=1.231e+07u
.ends

.subckt sky130_fd_pr__pfet_01v8_8DZSMJ a_n74_n100# a_16_n100# w_n212_n319# a_n33_n197#
X0 a_16_n100# a_n33_n197# a_n74_n100# w_n212_n319# sky130_fd_pr__pfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=160000u
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_D3C9B3 a_n36_n147# a_36_n50# w_n232_n269# a_n94_n50#
X0 a_36_n50# a_n36_n147# a_n94_n50# w_n232_n269# sky130_fd_pr__pfet_01v8_lvt ad=1.45e+11p pd=1.58e+06u as=1.45e+11p ps=1.58e+06u w=500000u l=360000u
.ends

.subckt vco ctrl out vcc gnd
Xsky130_fd_pr__nfet_01v8_Q8AFGD_1 m1_3250_1750# m1_970_1840# gnd gnd sky130_fd_pr__nfet_01v8_Q8AFGD
Xsky130_fd_pr__cap_mim_m3_1_9SN4GA_0 m1_3370_3860# gnd sky130_fd_pr__cap_mim_m3_1_9SN4GA
Xsky130_fd_pr__cap_mim_m3_1_9SN4GA_1 m1_970_3860# gnd sky130_fd_pr__cap_mim_m3_1_9SN4GA
Xx4 x4/A gnd vcc out gnd vcc sky130_fd_sc_hd__clkbuf_1
XXR40 vcc gnd m1_970_1840# sky130_fd_pr__res_xhigh_po_0p35_H4KU7R
XXM19 gnd m1_970_1840# m1_970_1840# gnd sky130_fd_pr__nfet_01v8_Q8AFGD
XXC30 m1_2570_3860# gnd sky130_fd_pr__cap_mim_m3_1_9SN4GA
XXR38 m1_n2285_5065# m1_970_1840# gnd sky130_fd_pr__res_xhigh_po_0p69_ET3NLF
XXM100 m1_2400_1760# m1_2570_3860# m1_3370_3860# gnd sky130_fd_pr__nfet_01v8_Q8AFGD
XXM102 m1_3145_3765# vcc vcc m1_970_4530# sky130_fd_pr__pfet_01v8_8DZSMJ
XXM105 m1_3250_1750# m1_3370_3860# x4/A gnd sky130_fd_pr__nfet_01v8_Q8AFGD
XXC29 m1_1770_3860# gnd sky130_fd_pr__cap_mim_m3_1_9SN4GA
XXM107 ctrl vcc vcc m1_n2285_5065# sky130_fd_pr__pfet_01v8_lvt_D3C9B3
XXM90 m1_850_1760# m1_970_3860# m1_1770_3860# gnd sky130_fd_pr__nfet_01v8_Q8AFGD
XXM91 m1_850_1760# m1_970_1840# gnd gnd sky130_fd_pr__nfet_01v8_Q8AFGD
XXM80 m1_970_4530# m1_970_1840# gnd gnd sky130_fd_pr__nfet_01v8_Q8AFGD
XXM92 m1_1525_3775# vcc vcc m1_970_4530# sky130_fd_pr__pfet_01v8_8DZSMJ
XXM82 m1_n75_3625# vcc vcc m1_970_4530# sky130_fd_pr__pfet_01v8_8DZSMJ
XXM81 vcc m1_970_4530# vcc m1_970_4530# sky130_fd_pr__pfet_01v8_8DZSMJ
XXM93 m1_1525_3775# m1_2570_3860# vcc m1_1770_3860# sky130_fd_pr__pfet_01v8_8DZSMJ
XXM83 m1_n75_3625# m1_970_3860# vcc x4/A sky130_fd_pr__pfet_01v8_8DZSMJ
XXM95 m1_1580_1770# m1_1770_3860# m1_2570_3860# gnd sky130_fd_pr__nfet_01v8_Q8AFGD
XXM96 m1_1580_1770# m1_970_1840# gnd gnd sky130_fd_pr__nfet_01v8_Q8AFGD
XXM85 m1_n60_1770# m1_970_1840# gnd gnd sky130_fd_pr__nfet_01v8_Q8AFGD
XXM97 m1_2375_3755# vcc vcc m1_970_4530# sky130_fd_pr__pfet_01v8_8DZSMJ
XXM86 m1_n60_1770# x4/A m1_970_3860# gnd sky130_fd_pr__nfet_01v8_Q8AFGD
XXM98 m1_2375_3755# m1_3370_3860# vcc m1_2570_3860# sky130_fd_pr__pfet_01v8_8DZSMJ
XXM87 m1_755_3765# vcc vcc m1_970_4530# sky130_fd_pr__pfet_01v8_8DZSMJ
Xsky130_fd_pr__pfet_01v8_8DZSMJ_0 m1_3145_3765# x4/A vcc m1_3370_3860# sky130_fd_pr__pfet_01v8_8DZSMJ
Xsky130_fd_pr__nfet_01v8_Q8AFGD_0 m1_2400_1760# m1_970_1840# gnd gnd sky130_fd_pr__nfet_01v8_Q8AFGD
XXM88 m1_755_3765# m1_1770_3860# vcc m1_970_3860# sky130_fd_pr__pfet_01v8_8DZSMJ
.ends

.subckt sky130_fd_pr__pfet_01v8_GXFJV8 a_n359_n2000# a_n301_n2097# w_n497_n2219# a_301_n2000#
X0 a_301_n2000# a_n301_n2097# a_n359_n2000# w_n497_n2219# sky130_fd_pr__pfet_01v8 ad=5.8e+12p pd=4.058e+07u as=5.8e+12p ps=4.058e+07u w=2e+07u l=3.01e+06u
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_2FRDLY c1_n1147_n1001# m3_n1187_n1041#
X0 c1_n1147_n1001# m3_n1187_n1041# sky130_fd_pr__cap_mim_m3_1 l=1.001e+07u w=1.001e+07u
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_XM7B29 a_n108_n1000# w_n246_n1219# a_n50_n1097#
+ a_50_n1000#
X0 a_50_n1000# a_n50_n1097# a_n108_n1000# w_n246_n1219# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+12p pd=2.058e+07u as=2.9e+12p ps=2.058e+07u w=1e+07u l=500000u
.ends

.subckt sky130_fd_pr__nfet_01v8_JFBZSQ a_n359_n2000# a_301_n2000# a_n461_n2174# a_n301_n2088#
X0 a_301_n2000# a_n301_n2088# a_n359_n2000# a_n461_n2174# sky130_fd_pr__nfet_01v8 ad=5.8e+12p pd=4.058e+07u as=5.8e+12p ps=4.058e+07u w=2e+07u l=3.01e+06u
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_XRYC29 a_n108_n1000# w_n246_n1219# a_n50_n1097#
+ a_50_n1000#
X0 a_50_n1000# a_n50_n1097# a_n108_n1000# w_n246_n1219# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+12p pd=2.058e+07u as=2.9e+12p ps=2.058e+07u w=1e+07u l=500000u
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_3LXTS5 a_n108_n300# w_n246_n519# a_n50_n397# a_50_n300#
X0 a_50_n300# a_n50_n397# a_n108_n300# w_n246_n519# sky130_fd_pr__pfet_01v8_lvt ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=500000u
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_ZSYV2F a_n35_3001# a_n165_n3563# a_n35_n3433#
X0 a_n35_n3433# a_n35_3001# a_n165_n3563# sky130_fd_pr__res_xhigh_po_0p35 l=3.001e+07u
.ends

.subckt user_analog_project_wrapper gpio_analog[0] gpio_analog[10] gpio_analog[11]
+ gpio_analog[12] gpio_analog[13] gpio_analog[14] gpio_analog[15] gpio_analog[16]
+ gpio_analog[17] gpio_analog[1] gpio_analog[2] gpio_analog[3] gpio_analog[4] gpio_analog[5]
+ gpio_analog[6] gpio_analog[7] gpio_analog[8] gpio_analog[9] gpio_noesd[0] gpio_noesd[10]
+ gpio_noesd[11] gpio_noesd[12] gpio_noesd[13] gpio_noesd[14] gpio_noesd[15] gpio_noesd[16]
+ gpio_noesd[17] gpio_noesd[1] gpio_noesd[2] gpio_noesd[3] gpio_noesd[4] gpio_noesd[5]
+ gpio_noesd[6] gpio_noesd[7] gpio_noesd[8] gpio_noesd[9] io_analog[0] io_analog[10]
+ io_analog[1] io_analog[2] io_analog[3] io_analog[7] io_analog[8] io_analog[9] io_analog[4]
+ io_analog[5] io_analog[6] io_clamp_high[0] io_clamp_high[1] io_clamp_high[2] io_clamp_low[0]
+ io_clamp_low[1] io_clamp_low[2] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_in_3v3[0] io_in_3v3[10] io_in_3v3[11] io_in_3v3[12]
+ io_in_3v3[13] io_in_3v3[14] io_in_3v3[15] io_in_3v3[16] io_in_3v3[17] io_in_3v3[18]
+ io_in_3v3[19] io_in_3v3[1] io_in_3v3[20] io_in_3v3[21] io_in_3v3[22] io_in_3v3[23]
+ io_in_3v3[24] io_in_3v3[25] io_in_3v3[26] io_in_3v3[2] io_in_3v3[3] io_in_3v3[4]
+ io_in_3v3[5] io_in_3v3[6] io_in_3v3[7] io_in_3v3[8] io_in_3v3[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100] la_data_in[101]
+ la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106]
+ la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111]
+ la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116]
+ la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121]
+ la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126]
+ la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16]
+ la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21]
+ la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27]
+ la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32]
+ la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38]
+ la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43]
+ la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49]
+ la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54]
+ la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5]
+ la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65]
+ la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70]
+ la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76]
+ la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81]
+ la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87]
+ la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92]
+ la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98]
+ la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2]
+ vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
Xsky130_fd_pr__cap_mim_m3_1_P68BUM_4 vssd1 vdda1 sky130_fd_pr__cap_mim_m3_1_P68BUM
Xsky130_fd_pr__cap_mim_m3_1_P68BUM_5 vssd1 vdda1 sky130_fd_pr__cap_mim_m3_1_P68BUM
Xanalogsub_0 vdda1 analogsub_0/Vplus gpio_analog[11] analogsub_0/Vminus gilbert_1/NB
+ filter_1/input vssd1 analogsub
Xsky130_fd_pr__res_xhigh_po_0p35_R9FY7S_1 vssd1 filter_1/pb vssd1 sky130_fd_pr__res_xhigh_po_0p35_R9FY7S
Xsky130_fd_pr__res_xhigh_po_0p35_R9FY7S_0 gilbert_1/NB vdda1 vssd1 sky130_fd_pr__res_xhigh_po_0p35_R9FY7S
Xsky130_fd_pr__cap_mim_m3_1_REKGFF_0 vssd1 vdda1 sky130_fd_pr__cap_mim_m3_1_REKGFF
Xanalogsub_1 vdda1 analogsub_1/Vplus gpio_analog[11] analogsub_1/Vminus gilbert_1/NB
+ filter_0/input vssd1 analogsub
Xsky130_fd_pr__cap_mim_m3_1_REKGFF_1 vssd1 vdda1 sky130_fd_pr__cap_mim_m3_1_REKGFF
Xanalogsub_2 vdda1 opamp_1/output gpio_analog[11] analogsub_2/Vminus gilbert_1/NB
+ analogsub_2/vout vssd1 analogsub
Xsky130_fd_pr__cap_mim_m3_1_REKGFF_2 vssd1 vdda1 sky130_fd_pr__cap_mim_m3_1_REKGFF
Xsky130_fd_pr__cap_mim_m3_1_5B6GLN_0 vdda1 vssd1 sky130_fd_pr__cap_mim_m3_1_5B6GLN
Xsky130_fd_pr__cap_mim_m3_1_REKGFF_4 vssd1 vdda1 sky130_fd_pr__cap_mim_m3_1_REKGFF
Xsky130_fd_pr__cap_mim_m3_1_REKGFF_3 vssd1 gpio_analog[11] sky130_fd_pr__cap_mim_m3_1_REKGFF
Xsky130_fd_pr__cap_mim_m3_1_REKGFF_5 vssd1 vdda1 sky130_fd_pr__cap_mim_m3_1_REKGFF
Xquadgen_0 io_in[15] gilbert_0/LO- gilbert_0/LO+ gilbert_1/LO+ gilbert_1/LO- vdda1
+ vssd1 vdda1 vssd1 quadgen
Xsky130_fd_pr__cap_mim_m3_1_REKGFF_6 vssd1 vdda1 sky130_fd_pr__cap_mim_m3_1_REKGFF
Xsky130_fd_pr__cap_mim_m3_1_REKGFF_7 vssd1 vdda1 sky130_fd_pr__cap_mim_m3_1_REKGFF
Xsky130_fd_pr__nfet_01v8_lvt_U9BGXT_0 gilbert_1/NB gilbert_1/NB vssd1 vssd1 sky130_fd_pr__nfet_01v8_lvt_U9BGXT
Xclkdiv_0 io_out[13] phasecmp_0/a vdda1 vdda1 clkdiv_0/x6/D clkdiv_0/x7/D vdda1 vdda1
+ clkdiv_0/x5/D vssd1 clkdiv
Xphasecmp_0 phasecmp_0/a io_in[10] gpio_analog[4] vdda1 vssd1 vssd1 vdda1 phasecmp
Xsky130_fd_pr__res_xhigh_po_0p35_LU79P3_1 opamp_1/inv opamp_0/inv vssd1 sky130_fd_pr__res_xhigh_po_0p35_LU79P3
Xsky130_fd_pr__res_xhigh_po_0p35_LU79P3_0 opamp_1/output opamp_1/inv vssd1 sky130_fd_pr__res_xhigh_po_0p35_LU79P3
Xsky130_fd_pr__cap_mim_m3_1_PUMBUM_0 li_35675_258517# gpio_analog[13] gpio_analog[13]
+ li_35675_258517# gpio_analog[13] li_35675_258517# li_35675_258517# gpio_analog[13]
+ sky130_fd_pr__cap_mim_m3_1_PUMBUM
Xsky130_fd_pr__cap_mim_m3_1_PUMBUM_2 m1_34962_259860# m4_64136_273264# m4_64136_273264#
+ m1_34962_259860# m4_64136_273264# m1_34962_259860# m1_34962_259860# m4_64136_273264#
+ sky130_fd_pr__cap_mim_m3_1_PUMBUM
Xsky130_fd_pr__nfet_01v8_lvt_JDBWNB_0 m1_34962_259860# vssd1 vssd1 li_35675_258517#
+ sky130_fd_pr__nfet_01v8_lvt_JDBWNB
Xsky130_fd_pr__cap_mim_m3_1_PUMBUM_1 vssd1 filter_1/pb filter_1/pb vssd1 filter_1/pb
+ vssd1 vssd1 filter_1/pb sky130_fd_pr__cap_mim_m3_1_PUMBUM
Xsky130_fd_pr__cap_mim_m3_1_R8KP6D_0 gpio_analog[12] gpio_analog[12] opamp_0/inv opamp_0/inv
+ sky130_fd_pr__cap_mim_m3_1_R8KP6D
Xsky130_fd_pr__cap_mim_m3_1_PUMBUM_3 m1_67449_275949# gilbert_1/RF+ gilbert_1/RF+
+ m1_67449_275949# gilbert_1/RF+ m1_67449_275949# m1_67449_275949# gilbert_1/RF+ sky130_fd_pr__cap_mim_m3_1_PUMBUM
Xsky130_fd_pr__res_xhigh_po_0p35_G3F5X4_0 m4_64136_273264# vssd1 gpio_analog[11] sky130_fd_pr__res_xhigh_po_0p35_G3F5X4
Xsky130_fd_pr__res_xhigh_po_0p35_G3F5X4_1 gilbert_1/RF+ vssd1 gpio_analog[11] sky130_fd_pr__res_xhigh_po_0p35_G3F5X4
Xsky130_fd_pr__res_xhigh_po_5p73_P7BAXV_0 gpio_analog[11] vssd1 vdda1 sky130_fd_pr__res_xhigh_po_5p73_P7BAXV
Xsky130_fd_pr__cap_mim_m3_1_PUMBUM_4 vssd1 gilbert_1/NB gilbert_1/NB vssd1 gilbert_1/NB
+ vssd1 vssd1 gilbert_1/NB sky130_fd_pr__cap_mim_m3_1_PUMBUM
Xsky130_fd_pr__res_xhigh_po_0p35_G3F5X4_2 analogsub_0/Vminus vssd1 gpio_analog[11]
+ sky130_fd_pr__res_xhigh_po_0p35_G3F5X4
Xsky130_fd_pr__res_xhigh_po_5p73_P7BAXV_1 vssd1 vssd1 gpio_analog[11] sky130_fd_pr__res_xhigh_po_5p73_P7BAXV
Xsky130_fd_pr__cap_mim_m3_1_PUMBUM_5 vssd1 gpio_analog[11] gpio_analog[11] vssd1 gpio_analog[11]
+ vssd1 vssd1 gpio_analog[11] sky130_fd_pr__cap_mim_m3_1_PUMBUM
Xsky130_fd_pr__pfet_01v8_lvt_TDASS5_0 m1_34962_259860# li_35675_258517# vssd1 vdda1
+ sky130_fd_pr__pfet_01v8_lvt_TDASS5
Xopamp_0 vdda1 opamp_0/inv opamp_0/noninv opamp_0/inv vssd1 opamp
Xsky130_fd_pr__cap_mim_m3_1_PUMBUM_6 gilbert_0/IF+ analogsub_1/Vminus analogsub_1/Vminus
+ gilbert_0/IF+ analogsub_1/Vminus gilbert_0/IF+ gilbert_0/IF+ analogsub_1/Vminus
+ sky130_fd_pr__cap_mim_m3_1_PUMBUM
Xfilter_0 vdda1 filter_0/input filter_0/out filter_1/pb vssd1 filter
Xsky130_fd_pr__res_xhigh_po_0p35_G3F5X4_3 analogsub_0/Vplus vssd1 gpio_analog[11]
+ sky130_fd_pr__res_xhigh_po_0p35_G3F5X4
Xsky130_fd_pr__pfet_01v8_lvt_TDASS5_1 li_35675_258517# li_35675_258517# m1_34962_259860#
+ vdda1 sky130_fd_pr__pfet_01v8_lvt_TDASS5
Xopamp_1 vdda1 opamp_1/inv gpio_analog[12] opamp_1/output vssd1 opamp
Xfilter_1 vdda1 filter_1/input filter_1/out filter_1/pb vssd1 filter
Xsky130_fd_pr__res_xhigh_po_0p35_G3F5X4_4 analogsub_1/Vminus vssd1 gpio_analog[11]
+ sky130_fd_pr__res_xhigh_po_0p35_G3F5X4
Xsky130_fd_pr__cap_mim_m3_1_PUMBUM_7 gilbert_0/IF- analogsub_1/Vplus analogsub_1/Vplus
+ gilbert_0/IF- analogsub_1/Vplus gilbert_0/IF- gilbert_0/IF- analogsub_1/Vplus sky130_fd_pr__cap_mim_m3_1_PUMBUM
Xopamp_2 vdda1 gpio_analog[10] opamp_2/noninv gpio_analog[9] vssd1 opamp
Xsky130_fd_sc_hd__clkbuf_16_0 gpio_analog[1] vssd1 vdda1 io_out[9] vssd1 vdda1 sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_pr__cap_mim_m3_1_PUMBUM_8 gilbert_1/IF- analogsub_0/Vplus analogsub_0/Vplus
+ gilbert_1/IF- analogsub_0/Vplus gilbert_1/IF- gilbert_1/IF- analogsub_0/Vplus sky130_fd_pr__cap_mim_m3_1_PUMBUM
Xsky130_fd_pr__res_xhigh_po_0p35_G3F5X4_5 analogsub_1/Vplus vssd1 gpio_analog[11]
+ sky130_fd_pr__res_xhigh_po_0p35_G3F5X4
Xsky130_fd_sc_hd__clkbuf_16_1 vco_0/out vssd1 vdda1 io_out[13] vssd1 vdda1 sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_pr__cap_mim_m3_1_PUMBUM_9 gilbert_1/IF+ analogsub_0/Vminus analogsub_0/Vminus
+ gilbert_1/IF+ analogsub_0/Vminus gilbert_1/IF+ gilbert_1/IF+ analogsub_0/Vminus
+ sky130_fd_pr__cap_mim_m3_1_PUMBUM
Xgilbert_0 vdda1 gilbert_0/LO+ gilbert_0/LO- gilbert_1/RF+ gpio_analog[11] gilbert_0/IF+
+ gilbert_0/IF- gilbert_1/NB filter_1/pb vssd1 gilbert
Xsky130_fd_pr__res_xhigh_po_0p35_G3F5X4_6 opamp_0/noninv vssd1 gpio_analog[11] sky130_fd_pr__res_xhigh_po_0p35_G3F5X4
Xsky130_fd_pr__pfet_01v8_lvt_TRXTS5_1 filter_1/pb vdda1 m1_34962_259860# vdda1 sky130_fd_pr__pfet_01v8_lvt_TRXTS5
Xgilbert_1 vdda1 gilbert_1/LO+ gilbert_1/LO- gilbert_1/RF+ gpio_analog[11] gilbert_1/IF+
+ gilbert_1/IF- gilbert_1/NB filter_1/pb vssd1 gilbert
Xsky130_fd_pr__res_xhigh_po_0p35_G3F5X4_7 analogsub_2/Vminus vssd1 gpio_analog[11]
+ sky130_fd_pr__res_xhigh_po_0p35_G3F5X4
Xsky130_fd_pr__cap_mim_m3_1_PUMBUM_10 analogsub_2/vout opamp_2/noninv opamp_2/noninv
+ analogsub_2/vout opamp_2/noninv analogsub_2/vout analogsub_2/vout opamp_2/noninv
+ sky130_fd_pr__cap_mim_m3_1_PUMBUM
Xvco_0 gpio_analog[5] vco_0/out vdda1 vssd1 vco
Xsky130_fd_pr__cap_mim_m3_1_PUMBUM_11 filter_1/out opamp_0/noninv opamp_0/noninv filter_1/out
+ opamp_0/noninv filter_1/out filter_1/out opamp_0/noninv sky130_fd_pr__cap_mim_m3_1_PUMBUM
Xsky130_fd_pr__pfet_01v8_GXFJV8_0 vdda1 gpio_analog[0] vdda1 gpio_analog[1] sky130_fd_pr__pfet_01v8_GXFJV8
Xsky130_fd_pr__cap_mim_m3_1_PUMBUM_12 filter_0/out analogsub_2/Vminus analogsub_2/Vminus
+ filter_0/out analogsub_2/Vminus filter_0/out filter_0/out analogsub_2/Vminus sky130_fd_pr__cap_mim_m3_1_PUMBUM
Xsky130_fd_pr__cap_mim_m3_1_2FRDLY_0 vdda1 vssd1 sky130_fd_pr__cap_mim_m3_1_2FRDLY
Xsky130_fd_pr__pfet_01v8_lvt_XM7B29_0 m1_67449_275949# vdda1 filter_1/pb vdda1 sky130_fd_pr__pfet_01v8_lvt_XM7B29
Xsky130_fd_pr__nfet_01v8_JFBZSQ_0 gpio_analog[1] vssd1 vssd1 gpio_analog[0] sky130_fd_pr__nfet_01v8_JFBZSQ
Xsky130_fd_pr__pfet_01v8_lvt_XRYC29_0 m1_67449_275949# vdda1 m4_64136_273264# vssd1
+ sky130_fd_pr__pfet_01v8_lvt_XRYC29
Xsky130_fd_pr__cap_mim_m3_1_P68BUM_0 vssd1 gpio_analog[11] sky130_fd_pr__cap_mim_m3_1_P68BUM
Xsky130_fd_pr__pfet_01v8_lvt_3LXTS5_0 filter_1/pb vdda1 filter_1/pb vdda1 sky130_fd_pr__pfet_01v8_lvt_3LXTS5
Xsky130_fd_pr__cap_mim_m3_1_P68BUM_1 vdda1 vssd1 sky130_fd_pr__cap_mim_m3_1_P68BUM
Xsky130_fd_pr__cap_mim_m3_1_P68BUM_2 vssd1 vdda1 sky130_fd_pr__cap_mim_m3_1_P68BUM
Xsky130_fd_pr__res_xhigh_po_0p35_ZSYV2F_0 opamp_2/noninv vssd1 gpio_analog[11] sky130_fd_pr__res_xhigh_po_0p35_ZSYV2F
Xsky130_fd_pr__cap_mim_m3_1_P68BUM_3 gpio_analog[11] vssd1 sky130_fd_pr__cap_mim_m3_1_P68BUM
R0 io_oeb[15] vdda1 sky130_fd_pr__res_generic_m3 w=560000u l=530000u
R1 vdda1 io_oeb[10] sky130_fd_pr__res_generic_m3 w=560000u l=620000u
R2 vssd1 io_oeb[9] sky130_fd_pr__res_generic_m3 w=560000u l=560000u
R3 vssd1 io_oeb[13] sky130_fd_pr__res_generic_m3 w=560000u l=770000u
.ends

