magic
tech sky130A
magscale 1 2
timestamp 1672355014
<< error_p >>
rect -131 1832 -130 1866
rect -35 -1832 -34 1832
rect 130 -1832 131 1866
<< pwell >>
rect -201 -1998 201 1998
<< psubdiff >>
rect -165 1928 -69 1962
rect 69 1928 165 1962
rect -165 1866 -130 1928
rect 130 1866 165 1928
rect -165 -1928 -130 -1866
rect 130 -1928 165 -1866
rect -165 -1962 -69 -1928
rect 69 -1962 165 -1928
<< psubdiffcont >>
rect -69 1928 69 1962
rect -165 -1866 -130 1866
rect 130 -1866 165 1866
rect -69 -1962 69 -1928
<< xpolycontact >>
rect -35 1400 35 1832
rect -35 -1832 35 -1400
<< xpolyres >>
rect -35 -1400 35 1400
<< locali >>
rect -165 1928 -69 1962
rect 69 1928 165 1962
rect -165 1866 -130 1928
rect 130 1866 165 1928
rect -165 -1928 -130 -1866
rect 130 -1928 165 -1866
rect -165 -1962 -69 -1928
rect 69 -1962 165 -1928
<< viali >>
rect -19 1417 19 1814
rect -18 1416 18 1417
rect -18 -1417 18 -1416
rect -19 -1814 19 -1417
<< metal1 >>
rect -25 1814 25 1826
rect -25 1417 -19 1814
rect 19 1417 25 1814
rect -25 1416 -18 1417
rect 18 1416 25 1417
rect -25 1405 25 1416
rect -24 1404 24 1405
rect -24 -1405 24 -1404
rect -25 -1416 25 -1405
rect -25 -1417 -18 -1416
rect 18 -1417 25 -1416
rect -25 -1814 -19 -1417
rect 19 -1814 25 -1417
rect -25 -1826 25 -1814
<< res0p35 >>
rect -37 -1402 37 1402
<< properties >>
string FIXED_BBOX -148 -1945 148 1945
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 14.0 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 81.075k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
