magic
tech sky130A
magscale 1 2
timestamp 1671573989
<< metal3 >>
rect -3086 9032 3086 9060
rect -3086 3208 3002 9032
rect 3066 3208 3086 9032
rect -3086 3180 3086 3208
rect -3086 2912 3086 2940
rect -3086 -2912 3002 2912
rect 3066 -2912 3086 2912
rect -3086 -2940 3086 -2912
rect -3086 -3208 3086 -3180
rect -3086 -9032 3002 -3208
rect 3066 -9032 3086 -3208
rect -3086 -9060 3086 -9032
<< via3 >>
rect 3002 3208 3066 9032
rect 3002 -2912 3066 2912
rect 3002 -9032 3066 -3208
<< mimcap >>
rect -3046 8980 2754 9020
rect -3046 3260 -3006 8980
rect 2714 3260 2754 8980
rect -3046 3220 2754 3260
rect -3046 2860 2754 2900
rect -3046 -2860 -3006 2860
rect 2714 -2860 2754 2860
rect -3046 -2900 2754 -2860
rect -3046 -3260 2754 -3220
rect -3046 -8980 -3006 -3260
rect 2714 -8980 2754 -3260
rect -3046 -9020 2754 -8980
<< mimcapcontact >>
rect -3006 3260 2714 8980
rect -3006 -2860 2714 2860
rect -3006 -8980 2714 -3260
<< metal4 >>
rect -198 8981 -94 9180
rect 2982 9032 3086 9180
rect -3007 8980 2715 8981
rect -3007 3260 -3006 8980
rect 2714 3260 2715 8980
rect -3007 3259 2715 3260
rect -198 2861 -94 3259
rect 2982 3208 3002 9032
rect 3066 3208 3086 9032
rect 2982 2912 3086 3208
rect -3007 2860 2715 2861
rect -3007 -2860 -3006 2860
rect 2714 -2860 2715 2860
rect -3007 -2861 2715 -2860
rect -198 -3259 -94 -2861
rect 2982 -2912 3002 2912
rect 3066 -2912 3086 2912
rect 2982 -3208 3086 -2912
rect -3007 -3260 2715 -3259
rect -3007 -8980 -3006 -3260
rect 2714 -8980 2715 -3260
rect -3007 -8981 2715 -8980
rect -198 -9180 -94 -8981
rect 2982 -9032 3002 -3208
rect 3066 -9032 3086 -3208
rect 2982 -9180 3086 -9032
<< properties >>
string FIXED_BBOX -3086 3180 2794 9060
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 29.0 l 29.0 val 1.704k carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
