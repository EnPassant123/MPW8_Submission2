magic
tech sky130A
magscale 1 2
timestamp 1639841760
<< error_p >>
rect 5036 7870 5051 7898
rect 5008 7676 5023 7870
rect 20366 7862 20381 7890
rect 20394 7668 20409 7862
use example_por  example_por_0
timestamp 1639841760
transform -1 0 11285 0 1 -14
box 0 0 11344 8338
use example_por  example_por_1
timestamp 1639841760
transform 1 0 14132 0 1 -22
box 0 0 11344 8338
<< end >>
