magic
tech sky130A
timestamp 1671518644
<< metal3 >>
rect -793 706 793 720
rect -793 -706 751 706
rect 783 -706 793 706
rect -793 -720 793 -706
<< via3 >>
rect 751 -706 783 706
<< mimcap >>
rect -773 680 627 700
rect -773 -680 -753 680
rect 607 -680 627 680
rect -773 -700 627 -680
<< mimcapcontact >>
rect -753 -680 607 680
<< metal4 >>
rect 743 706 791 714
rect 743 -706 751 706
rect 783 -706 791 706
rect 743 -714 791 -706
<< properties >>
string FIXED_BBOX -793 -720 647 720
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 14.0 l 14.0 val 402.64 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
