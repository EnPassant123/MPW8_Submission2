magic
tech sky130A
magscale 1 2
timestamp 1672366774
<< nwell >>
rect -109 -691 790 -370
rect 2471 -691 3420 -370
rect 4430 -691 5080 -370
rect -109 -770 212 -691
rect -1860 -806 212 -770
rect -1900 -1091 212 -806
rect 4759 -1140 5080 -691
rect 4499 -1370 5080 -1140
rect 2471 -1691 3630 -1370
rect 4335 -1461 5080 -1370
rect 4335 -1691 4820 -1461
<< pwell >>
rect 319 -971 781 -789
rect 2560 -931 3451 -749
rect 319 -1149 501 -971
rect -1861 -1331 501 -1149
rect 319 -1799 501 -1331
rect 319 -1981 711 -1799
rect 2560 -1931 3471 -1749
<< locali >>
rect 4589 -403 4804 -391
rect 4587 -438 4804 -403
rect 389 -621 577 -551
rect 507 -633 577 -621
rect 4769 -611 4804 -438
rect 4769 -621 5049 -611
rect 507 -703 726 -633
rect 4769 -650 5056 -621
rect 2686 -737 3326 -697
rect 351 -927 385 -799
rect 4525 -805 4664 -729
rect -1008 -953 -824 -946
rect -1008 -1006 -884 -953
rect -831 -1006 -824 -953
rect 123 -961 385 -927
rect -1008 -1011 -824 -1006
rect -1008 -1094 -943 -1011
rect 5177 -1043 7294 -1037
rect 5177 -1081 7250 -1043
rect 7288 -1081 7294 -1043
rect 5177 -1087 7294 -1081
rect -1412 -1097 -1276 -1096
rect -1545 -1103 -1276 -1097
rect -1545 -1157 -1539 -1103
rect -1485 -1141 -1276 -1103
rect -1174 -1136 -943 -1094
rect -1008 -1138 -943 -1136
rect -808 -1137 -505 -1097
rect -1485 -1157 -1407 -1141
rect -1545 -1163 -1407 -1157
rect -808 -1218 -768 -1137
rect -1118 -1258 -768 -1218
rect 129 -1281 293 -1247
rect 259 -1523 293 -1281
rect 179 -1557 293 -1523
rect 179 -1765 213 -1557
rect 5179 -1511 7304 -1505
rect 5179 -1553 7256 -1511
rect 7298 -1553 7304 -1511
rect 5179 -1559 7304 -1553
rect 409 -1703 726 -1633
rect 2706 -1737 2726 -1697
rect 2994 -1737 3326 -1697
rect 931 -1799 957 -1765
rect 2994 -2046 3034 -1737
rect 4525 -1805 4732 -1729
rect 4589 -1940 5044 -1935
rect 4589 -1969 5096 -1940
rect 7359 -1964 7670 -1922
<< viali >>
rect 2373 -747 2439 -681
rect 351 -799 385 -765
rect 939 -799 973 -765
rect 4664 -805 4740 -729
rect -884 -1006 -831 -953
rect 5127 -1087 5177 -1037
rect 7250 -1081 7288 -1043
rect -1539 -1157 -1485 -1103
rect 5125 -1559 5179 -1505
rect 7256 -1553 7298 -1511
rect 2373 -1745 2439 -1679
rect 179 -1799 213 -1765
rect 957 -1799 991 -1765
rect 4732 -1805 4808 -1729
rect 2994 -2086 3034 -2046
<< metal1 >>
rect 157 -395 655 -359
rect 157 -453 759 -395
rect 2721 -418 3451 -360
rect 157 -601 215 -453
rect 2733 -456 3359 -418
rect 4612 -456 5354 -360
rect 151 -659 157 -601
rect 215 -659 221 -601
rect -1818 -818 -349 -760
rect 157 -798 215 -659
rect 5216 -668 5312 -456
rect 2361 -681 2451 -675
rect 2361 -687 2373 -681
rect 2439 -687 2451 -681
rect 2361 -753 2367 -687
rect 2445 -753 2451 -687
rect 4658 -729 4746 -717
rect 2367 -759 2445 -753
rect -1818 -856 -441 -818
rect 53 -856 215 -798
rect 339 -765 397 -759
rect 339 -799 351 -765
rect 385 -768 397 -765
rect 927 -765 985 -759
rect 927 -768 939 -765
rect 385 -796 939 -768
rect 385 -799 397 -796
rect 339 -805 397 -799
rect 927 -799 939 -796
rect 973 -768 985 -765
rect 973 -796 1594 -768
rect 973 -799 985 -796
rect 927 -805 985 -799
rect 4658 -805 4664 -729
rect 4740 -799 5174 -729
rect 5216 -764 7200 -668
rect 4740 -805 5177 -799
rect 4658 -817 4746 -805
rect -896 -1012 -890 -947
rect -825 -1012 -819 -947
rect 349 -1000 759 -911
rect 2731 -942 3359 -904
rect 2689 -1000 3451 -942
rect -1545 -1097 -1479 -1091
rect -1551 -1163 -1545 -1097
rect -1479 -1163 -1473 -1097
rect -1545 -1169 -1479 -1163
rect -1794 -1354 -1346 -1306
rect -1119 -1342 -441 -1309
rect -1794 -1369 -1332 -1354
rect -1816 -1400 -1285 -1369
rect -1131 -1400 -441 -1342
rect 349 -1351 407 -1000
rect 5127 -1025 5177 -805
rect 5220 -910 7200 -814
rect 7250 -880 7294 -754
rect 5121 -1037 5183 -1025
rect 5121 -1087 5127 -1037
rect 5177 -1087 5183 -1037
rect 5121 -1099 5183 -1087
rect -119 -1381 -61 -1361
rect -119 -1907 -33 -1381
rect 63 -1409 407 -1351
rect 497 -1418 503 -1360
rect 561 -1418 759 -1360
rect 2683 -1418 3359 -1360
rect 2697 -1456 3359 -1418
rect 5119 -1505 5185 -1493
rect 5119 -1559 5125 -1505
rect 5179 -1559 5185 -1505
rect 5119 -1571 5185 -1559
rect 2361 -1679 2451 -1673
rect 2361 -1685 2373 -1679
rect 2439 -1685 2451 -1679
rect 2361 -1751 2367 -1685
rect 2445 -1751 2451 -1685
rect 4726 -1729 4814 -1717
rect 5125 -1729 5179 -1571
rect 173 -1765 219 -1753
rect 2367 -1757 2445 -1751
rect 173 -1799 179 -1765
rect 213 -1768 219 -1765
rect 945 -1765 1003 -1759
rect 945 -1768 957 -1765
rect 213 -1796 957 -1768
rect 213 -1799 219 -1796
rect 173 -1811 219 -1799
rect 945 -1799 957 -1796
rect 991 -1768 1003 -1765
rect 991 -1796 1570 -1768
rect 991 -1799 1003 -1796
rect 945 -1805 1003 -1799
rect 4726 -1805 4732 -1729
rect 4808 -1783 5179 -1729
rect 5232 -1666 5328 -910
rect 7104 -1216 7200 -910
rect 7244 -1043 7294 -880
rect 7244 -1081 7250 -1043
rect 7288 -1081 7294 -1043
rect 7244 -1093 7294 -1081
rect 7104 -1312 7960 -1216
rect 7104 -1666 7200 -1312
rect 5232 -1668 7200 -1666
rect 7250 -1511 7304 -1499
rect 7250 -1553 7256 -1511
rect 7298 -1553 7304 -1511
rect 5232 -1764 7208 -1668
rect 4808 -1805 5172 -1783
rect 4726 -1817 4814 -1805
rect -119 -2000 759 -1907
rect 2697 -1942 3359 -1905
rect 4606 -1907 4682 -1904
rect 5221 -1907 7210 -1814
rect 7250 -1858 7304 -1553
rect 9228 -1844 9838 -686
rect 2633 -2000 3379 -1942
rect 4589 -2000 5396 -1907
rect 2988 -2040 3040 -2034
rect 2982 -2092 2988 -2040
rect 3040 -2092 3046 -2040
rect 2988 -2098 3040 -2092
<< via1 >>
rect 157 -659 215 -601
rect 2367 -747 2373 -687
rect 2373 -747 2439 -687
rect 2439 -747 2445 -687
rect 2367 -753 2445 -747
rect -890 -953 -825 -947
rect -890 -1006 -884 -953
rect -884 -1006 -831 -953
rect -831 -1006 -825 -953
rect -890 -1012 -825 -1006
rect -1545 -1103 -1479 -1097
rect -1545 -1157 -1539 -1103
rect -1539 -1157 -1485 -1103
rect -1485 -1157 -1479 -1103
rect -1545 -1163 -1479 -1157
rect 503 -1418 561 -1360
rect 2367 -1745 2373 -1685
rect 2373 -1745 2439 -1685
rect 2439 -1745 2445 -1685
rect 2367 -1751 2445 -1745
rect 2988 -2046 3040 -2040
rect 2988 -2086 2994 -2046
rect 2994 -2086 3034 -2046
rect 3034 -2086 3040 -2046
rect 2988 -2092 3040 -2086
<< metal2 >>
rect -890 -306 2439 -241
rect -890 -947 -825 -306
rect 157 -601 215 -595
rect 157 -925 215 -659
rect 2373 -687 2439 -306
rect 2361 -753 2367 -687
rect 2445 -753 2451 -687
rect 157 -983 561 -925
rect -890 -1018 -825 -1012
rect -1551 -1163 -1545 -1097
rect -1479 -1163 -1473 -1097
rect -1545 -2097 -1479 -1163
rect 503 -1360 561 -983
rect 503 -1424 561 -1418
rect 2361 -1751 2367 -1685
rect 2445 -1751 2451 -1685
rect 2373 -2046 2439 -1751
rect 2988 -2040 3040 -2034
rect 2373 -2086 2988 -2046
rect 2373 -2097 2439 -2086
rect -1545 -2163 2439 -2097
rect 2988 -2098 3040 -2092
use sky130_fd_pr__pfet_01v8_QP79FH  XM108
timestamp 1672366774
transform 0 -1 6219 1 0 -787
box -212 -1219 212 1219
use sky130_fd_pr__nfet_01v8_A5ES5P  XM109
timestamp 1672366774
transform 0 1 6210 -1 0 -1789
box -211 -1210 211 1210
use sky130_fd_pr__res_xhigh_po_5p73_WAQYE6  XR17
timestamp 1672366774
transform 0 1 8714 -1 0 -1261
box -739 -1114 739 1114
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1672366774
transform 1 0 -1862 0 1 -1352
box -38 -48 130 592
use sky130_fd_sc_hd__dfrbp_1  x28 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1672366774
transform 1 0 638 0 1 -1952
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrbp_1  x29
timestamp 1672366774
transform 1 0 638 0 1 -952
box -38 -48 2154 592
use sky130_fd_sc_hd__bufbuf_8  x30 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1672366774
transform 1 0 3238 0 1 -1952
box -38 -48 1418 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  x31 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1672366774
transform 1 0 -562 0 1 -1352
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  x39 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1672366774
transform 1 0 -1362 0 1 -1352
box -38 -48 314 592
use sky130_fd_sc_hd__bufbuf_8  x162
timestamp 1672366774
transform 1 0 3238 0 1 -952
box -38 -48 1418 592
<< labels >>
rlabel metal1 5120 -434 5152 -404 1 vcc
port 0 n
rlabel locali 412 -604 444 -574 1 a
port 1 n
rlabel locali 448 -1682 480 -1652 1 b
port 2 n
rlabel metal1 9698 -1644 9730 -1614 1 out
port 3 n
rlabel locali 7512 -1956 7524 -1942 1 ground
port 4 n
<< end >>
