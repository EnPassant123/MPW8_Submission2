magic
tech sky130A
magscale 1 2
timestamp 1672366615
<< nwell >>
rect -247 -519 247 519
<< pmoslvt >>
rect -51 -300 51 300
<< pdiff >>
rect -109 288 -51 300
rect -109 -288 -97 288
rect -63 -288 -51 288
rect -109 -300 -51 -288
rect 51 288 109 300
rect 51 -288 63 288
rect 97 -288 109 288
rect 51 -300 109 -288
<< pdiffc >>
rect -97 -288 -63 288
rect 63 -288 97 288
<< nsubdiff >>
rect -211 449 -115 483
rect 115 449 211 483
rect -211 387 -177 449
rect 177 387 211 449
rect -211 -449 -177 -387
rect 177 -449 211 -387
rect -211 -483 -115 -449
rect 115 -483 211 -449
<< nsubdiffcont >>
rect -115 449 115 483
rect -211 -387 -177 387
rect 177 -387 211 387
rect -115 -483 115 -449
<< poly >>
rect -51 381 51 397
rect -51 347 -35 381
rect 35 347 51 381
rect -51 300 51 347
rect -51 -347 51 -300
rect -51 -381 -35 -347
rect 35 -381 51 -347
rect -51 -397 51 -381
<< polycont >>
rect -35 347 35 381
rect -35 -381 35 -347
<< locali >>
rect -211 449 -115 483
rect 115 449 211 483
rect -211 387 -177 449
rect 177 387 211 449
rect -51 347 -35 381
rect 35 347 51 381
rect -97 288 -63 304
rect -97 -304 -63 -288
rect 63 288 97 304
rect 63 -304 97 -288
rect -51 -381 -35 -347
rect 35 -381 51 -347
rect -211 -449 -177 -387
rect 177 -449 211 -387
rect -211 -483 -115 -449
rect 115 -483 211 -449
<< viali >>
rect -35 347 35 381
rect -97 -288 -63 288
rect 63 -288 97 288
rect -35 -381 35 -347
<< metal1 >>
rect -47 381 47 387
rect -47 347 -35 381
rect 35 347 47 381
rect -47 341 47 347
rect -103 288 -57 300
rect -103 -288 -97 288
rect -63 -288 -57 288
rect -103 -300 -57 -288
rect 57 288 103 300
rect 57 -288 63 288
rect 97 -288 103 288
rect 57 -300 103 -288
rect -47 -347 47 -341
rect -47 -381 -35 -347
rect 35 -381 47 -347
rect -47 -387 47 -381
<< properties >>
string FIXED_BBOX -194 -466 194 466
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 3.0 l 0.505 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
