magic
tech sky130A
magscale 1 2
timestamp 1672367450
<< nwell >>
rect 3951 3010 4754 3331
<< pwell >>
rect 4077 3415 4716 3571
<< locali >>
rect -1815 5735 -1415 5785
rect -2155 5715 -1415 5735
rect -2155 5665 -1745 5715
rect -1485 5709 -1415 5715
rect -1485 5651 -1479 5709
rect -1421 5651 -1415 5709
rect -1485 5645 -1415 5651
rect -1640 5374 -1580 5560
rect -1640 5326 -1634 5374
rect -1586 5326 -1580 5374
rect -1640 5320 -1580 5326
rect 570 5157 610 5160
rect 570 5123 573 5157
rect 607 5123 610 5157
rect 570 5020 610 5123
rect 1370 5157 1410 5160
rect 1370 5123 1373 5157
rect 1407 5123 1410 5157
rect 1370 5020 1410 5123
rect 2150 5157 2190 5160
rect 2150 5123 2153 5157
rect 2187 5123 2190 5157
rect 2150 5020 2190 5123
rect 2860 5020 2900 5110
rect -690 4980 3500 5020
rect -220 4010 -180 4980
rect 570 4800 610 4980
rect 1370 4810 1410 4980
rect 2150 4810 2190 4980
rect 2860 4820 2900 4980
rect -220 3970 3520 4010
rect 3670 3377 4030 3380
rect 3670 3343 3673 3377
rect 3707 3343 4030 3377
rect 4183 3353 4357 3387
rect 3670 3340 4030 3343
rect 230 3267 3710 3270
rect 230 3233 3673 3267
rect 3707 3233 3710 3267
rect 230 3230 3710 3233
rect 130 2440 3490 2480
rect -1570 2230 -1090 2270
rect -1570 1480 -1530 2230
rect -1145 2119 -610 2125
rect -1145 2081 -654 2119
rect -616 2081 -610 2119
rect -1145 2075 -610 2081
rect -306 1657 -266 1660
rect -306 1623 -303 1657
rect -269 1623 -266 1657
rect -306 1480 -266 1623
rect 490 1480 530 1620
rect 640 1480 680 2440
rect 1300 1480 1340 1630
rect 2040 1480 2080 1620
rect 2870 1480 2910 1630
rect -2170 1440 3580 1480
rect -434 1410 -340 1440
rect -380 1337 -340 1410
rect -380 1303 -377 1337
rect -343 1303 -340 1337
rect -380 1300 -340 1303
rect 490 1337 530 1440
rect 490 1303 493 1337
rect 527 1303 530 1337
rect 490 1300 530 1303
rect 1300 1337 1340 1440
rect 1300 1303 1303 1337
rect 1337 1303 1340 1337
rect 1300 1300 1340 1303
rect 2040 1337 2080 1440
rect 2040 1303 2043 1337
rect 2077 1303 2080 1337
rect 2040 1300 2080 1303
rect 2870 1337 2910 1440
rect 2870 1303 2873 1337
rect 2907 1303 2910 1337
rect 2870 1300 2910 1303
<< viali >>
rect -1479 5651 -1421 5709
rect -1640 5560 -1580 5620
rect -1634 5326 -1586 5374
rect 573 5123 607 5157
rect 1373 5123 1407 5157
rect 2153 5123 2187 5157
rect 2860 5110 2900 5150
rect 570 4760 610 4800
rect 1370 4770 1410 4810
rect 2150 4770 2190 4810
rect 2860 4780 2900 4820
rect 3673 3343 3707 3377
rect 190 3230 230 3270
rect 3673 3233 3707 3267
rect -1195 2075 -1145 2125
rect -654 2081 -616 2119
rect -303 1623 -269 1657
rect 490 1620 530 1660
rect 1300 1630 1340 1670
rect 2040 1620 2080 1660
rect 2870 1630 2910 1670
rect -377 1303 -343 1337
rect 493 1303 527 1337
rect 1303 1303 1337 1337
rect 2043 1303 2077 1337
rect 2873 1303 2907 1337
<< metal1 >>
rect -1260 6080 -720 6220
rect -1260 5715 -1120 6080
rect -1525 5709 -1120 5715
rect -1525 5651 -1479 5709
rect -1421 5651 -1120 5709
rect -1525 5645 -1120 5651
rect -1652 5620 -1568 5626
rect -2000 5560 -1640 5620
rect -1580 5560 -1568 5620
rect -1652 5554 -1568 5560
rect -1525 5510 -1455 5645
rect -1260 5560 -1120 5645
rect -2080 5505 -2010 5510
rect -2285 5435 -2010 5505
rect -2285 5135 -2215 5435
rect -2080 5420 -2010 5435
rect -1920 5440 -1455 5510
rect -1920 5420 -1850 5440
rect -1640 5380 -1580 5386
rect -2020 5374 -1580 5380
rect -2020 5326 -1634 5374
rect -1586 5326 -1580 5374
rect -2020 5320 -1580 5326
rect -1640 5314 -1580 5320
rect -860 5260 -720 6080
rect -880 5250 3640 5260
rect -880 5190 3880 5250
rect -880 5157 3640 5190
rect -2285 5065 -1865 5135
rect -880 5123 573 5157
rect 607 5123 1373 5157
rect 1407 5123 2153 5157
rect 2187 5150 3640 5157
rect 2187 5123 2860 5150
rect -880 5110 2860 5123
rect 2900 5110 3640 5150
rect -2050 4450 -1870 5065
rect -880 4670 -840 5110
rect 2848 5104 2912 5110
rect 3500 5030 3540 5110
rect 3500 4990 3620 5030
rect -660 4860 3440 4900
rect -650 4670 -610 4810
rect -880 4630 -610 4670
rect -570 4575 -530 4860
rect 135 4665 185 4815
rect -615 4570 -530 4575
rect -620 4530 -530 4570
rect -75 4615 185 4665
rect 240 4800 280 4810
rect 564 4800 616 4812
rect 240 4760 570 4800
rect 610 4760 616 4800
rect 240 4630 280 4760
rect 564 4748 616 4760
rect 935 4665 985 4815
rect 1364 4810 1416 4822
rect 2854 4820 2906 4832
rect 3580 4820 3620 4990
rect 755 4615 985 4665
rect 1030 4770 1370 4810
rect 1410 4770 1416 4810
rect 1030 4620 1070 4770
rect 1364 4758 1416 4770
rect 1735 4665 1785 4815
rect 2138 4810 2202 4816
rect 1525 4615 1785 4665
rect 1840 4770 2150 4810
rect 2190 4770 2202 4810
rect 1840 4620 1880 4770
rect 2138 4764 2202 4770
rect 2545 4675 2595 4815
rect 2375 4625 2595 4675
rect 2640 4780 2860 4820
rect 2900 4780 2906 4820
rect 2640 4630 2680 4780
rect 2854 4768 2906 4780
rect 3335 4665 3385 4805
rect -1250 2260 -1160 2800
rect -615 2295 -565 4530
rect -75 3675 -25 4615
rect 170 4530 260 4580
rect 170 3860 260 3900
rect 755 3815 805 4615
rect 970 4530 1060 4580
rect 970 3860 1060 3900
rect 1525 3825 1575 4615
rect 1770 4530 1860 4580
rect 1770 3860 1860 3900
rect 135 3675 185 3815
rect -75 3670 185 3675
rect 230 3670 270 3810
rect 755 3765 985 3815
rect -75 3625 190 3670
rect 230 3630 560 3670
rect 100 3620 190 3625
rect 520 3580 560 3630
rect 935 3625 985 3765
rect 1040 3660 1080 3820
rect 1525 3775 1785 3825
rect 1040 3620 1380 3660
rect 1340 3580 1380 3620
rect 1735 3615 1785 3775
rect 1830 3670 1870 3810
rect 2375 3805 2425 4625
rect 3145 4615 3385 4665
rect 3430 4780 3620 4820
rect 3430 4630 3470 4780
rect 2570 4530 2660 4580
rect 2570 3860 2660 3900
rect 3145 3815 3195 4615
rect 3370 4530 3460 4580
rect 3370 3860 3460 3900
rect 2375 3755 2585 3805
rect 1830 3630 2150 3670
rect 190 3276 230 3570
rect 520 3540 1040 3580
rect 1340 3540 1840 3580
rect 2110 3560 2150 3630
rect 2535 3625 2585 3755
rect 2640 3660 2680 3810
rect 3145 3765 3395 3815
rect 2640 3620 3040 3660
rect 3000 3570 3040 3620
rect 3345 3615 3395 3765
rect 3430 3660 3470 3810
rect 3820 3766 3880 5190
rect 3820 3706 4820 3766
rect 3430 3620 3710 3660
rect 178 3270 242 3276
rect 178 3230 190 3270
rect 230 3230 242 3270
rect 178 3224 242 3230
rect 190 2840 230 3224
rect 520 2890 560 3540
rect 520 2850 1040 2890
rect 1340 2880 1380 3540
rect 2110 3520 2640 3560
rect 3000 3530 3450 3570
rect 2110 2890 2150 3520
rect 3000 2890 3040 3530
rect 3670 3383 3710 3620
rect 3661 3377 3719 3383
rect 3661 3343 3673 3377
rect 3707 3343 3719 3377
rect 3661 3337 3719 3343
rect 3670 3273 3710 3337
rect 3667 3267 3713 3273
rect 3667 3233 3673 3267
rect 3707 3233 3713 3267
rect 3667 3227 3713 3233
rect 140 2660 190 2810
rect -1505 2170 -1160 2260
rect -915 2245 -565 2295
rect -60 2620 190 2660
rect 230 2660 280 2800
rect 520 2672 560 2850
rect 1340 2840 1840 2880
rect 2110 2850 2650 2890
rect 3000 2850 3470 2890
rect 494 2666 560 2672
rect 230 2620 494 2660
rect -1505 2075 -1415 2170
rect -1207 2125 -1133 2131
rect -1207 2075 -1195 2125
rect -1145 2075 -1133 2125
rect -1505 2069 -1133 2075
rect -1505 2025 -1145 2069
rect -2040 1595 -1870 2010
rect -1505 1595 -1415 2025
rect -1195 1905 -1145 2025
rect -1195 1855 -1115 1905
rect -1250 1650 -1210 1800
rect -2040 1510 -1415 1595
rect -1955 1505 -1415 1510
rect -1360 1610 -1210 1650
rect -1360 1350 -1320 1610
rect -1165 1535 -1115 1855
rect -915 1670 -865 2245
rect -660 2119 -610 2131
rect -660 2081 -654 2119
rect -616 2081 -610 2119
rect -660 1890 -610 2081
rect -660 1840 -530 1890
rect -60 1810 -20 2620
rect 230 2610 280 2620
rect 546 2620 560 2666
rect 950 2650 990 2800
rect 1340 2692 1380 2840
rect 1334 2686 1386 2692
rect 494 2608 546 2614
rect 850 2610 990 2650
rect 1030 2634 1334 2660
rect 1750 2650 1790 2800
rect 1030 2628 1386 2634
rect 1030 2620 1380 2628
rect 1580 2610 1790 2650
rect 1830 2660 1870 2810
rect 2110 2692 2150 2850
rect 2104 2686 2156 2692
rect 1830 2634 2104 2660
rect 2550 2660 2590 2800
rect 2640 2660 2680 2800
rect 3000 2672 3040 2850
rect 2994 2666 3046 2672
rect 1830 2628 2156 2634
rect 1830 2620 2150 2628
rect 2400 2620 2590 2660
rect 2630 2620 2994 2660
rect 170 2530 260 2570
rect 170 1840 260 1890
rect -665 1670 -615 1805
rect -915 1620 -610 1670
rect -570 1660 -530 1800
rect -60 1770 190 1810
rect -315 1660 -257 1663
rect -570 1657 -257 1660
rect -570 1623 -303 1657
rect -269 1623 -257 1657
rect -570 1620 -257 1623
rect -315 1617 -257 1620
rect 150 1610 190 1770
rect 240 1660 280 1810
rect 850 1800 890 2610
rect 960 2530 1050 2570
rect 970 1840 1060 1890
rect 1580 1810 1620 2610
rect 1760 2530 1850 2570
rect 1770 1840 1860 1890
rect 850 1760 990 1800
rect 478 1660 542 1666
rect 240 1620 490 1660
rect 530 1620 542 1660
rect 950 1620 990 1760
rect 1040 1670 1080 1810
rect 1580 1770 1790 1810
rect 2400 1800 2440 2620
rect 3350 2650 3390 2810
rect 3440 2660 3480 2800
rect 3670 2660 3710 3227
rect 3820 3060 3880 3706
rect 4626 3640 4686 3644
rect 4113 3584 4686 3640
rect 4113 3582 4663 3584
rect 4341 3071 4399 3582
rect 4760 3072 4820 3706
rect 4626 3071 4820 3072
rect 3820 3000 4020 3060
rect 4341 3013 4406 3071
rect 4586 3013 4820 3071
rect 2994 2608 3046 2614
rect 3250 2610 3390 2650
rect 3430 2620 3710 2660
rect 2570 2540 2660 2580
rect 2560 1840 2650 1890
rect 1288 1670 1352 1676
rect 1040 1630 1300 1670
rect 1340 1630 1352 1670
rect 478 1614 542 1620
rect 1040 1610 1080 1630
rect 1288 1624 1352 1630
rect 1750 1620 1790 1770
rect 1840 1660 1880 1800
rect 2400 1760 2590 1800
rect 2028 1660 2092 1666
rect 1840 1620 2040 1660
rect 2080 1620 2092 1660
rect 2550 1620 2590 1760
rect 2630 1670 2670 1810
rect 3250 1790 3290 2610
rect 3370 2540 3460 2580
rect 3370 1840 3460 1890
rect 3335 1790 3386 1796
rect 3250 1750 3386 1790
rect 2858 1670 2922 1676
rect 2630 1630 2870 1670
rect 2910 1630 2922 1670
rect 2630 1620 2670 1630
rect 2858 1624 2922 1630
rect 2028 1614 2092 1620
rect 3335 1615 3386 1750
rect 3430 1660 3470 1800
rect 3430 1620 3690 1660
rect -650 1530 3450 1570
rect 2995 1350 3145 1356
rect 3650 1350 3690 1620
rect -1400 1337 655 1350
rect -1400 1310 -377 1337
rect -390 1303 -377 1310
rect -343 1303 493 1337
rect 527 1303 655 1337
rect -390 1200 655 1303
rect 805 1337 2995 1350
rect 805 1303 1303 1337
rect 1337 1303 2043 1337
rect 2077 1303 2873 1337
rect 2907 1303 2995 1337
rect 805 1200 2995 1303
rect 3145 1349 4130 1350
rect 4341 1349 4399 3013
rect 4626 3012 4820 3013
rect 3145 1291 4399 1349
rect 3145 1200 4130 1291
rect 630 1190 670 1200
rect 2995 1194 3145 1200
<< via1 >>
rect 494 2614 546 2666
rect 1334 2634 1386 2686
rect 2104 2634 2156 2686
rect 2994 2614 3046 2666
rect 655 1200 805 1350
rect 2995 1200 3145 1350
<< metal2 >>
rect 1330 2690 1390 2699
rect 2100 2690 2160 2699
rect 490 2670 550 2679
rect 488 2614 490 2666
rect 550 2614 552 2666
rect 1328 2634 1330 2686
rect 1390 2634 1392 2686
rect 2098 2634 2100 2686
rect 2160 2634 2162 2686
rect 2990 2670 3050 2679
rect 1330 2621 1390 2630
rect 2100 2621 2160 2630
rect 2988 2614 2990 2666
rect 3050 2614 3052 2666
rect 490 2601 550 2610
rect 2990 2601 3050 2610
rect 2981 1430 2990 1490
rect 3050 1430 3370 1490
rect 655 1350 805 1359
rect 2995 1350 3145 1359
rect 2989 1200 2995 1350
rect 3145 1200 3151 1350
rect 655 1191 805 1200
rect 2995 1191 3145 1200
rect 3310 1178 3370 1430
rect 3310 1122 3312 1178
rect 3368 1122 3370 1178
rect 3310 1120 3370 1122
rect 3312 1113 3368 1120
<< via2 >>
rect 1330 2686 1390 2690
rect 2100 2686 2160 2690
rect 490 2666 550 2670
rect 490 2614 494 2666
rect 494 2614 546 2666
rect 546 2614 550 2666
rect 1330 2634 1334 2686
rect 1334 2634 1386 2686
rect 1386 2634 1390 2686
rect 2100 2634 2104 2686
rect 2104 2634 2156 2686
rect 2156 2634 2160 2686
rect 2990 2666 3050 2670
rect 1330 2630 1390 2634
rect 2100 2630 2160 2634
rect 2990 2614 2994 2666
rect 2994 2614 3046 2666
rect 3046 2614 3050 2666
rect 490 2610 550 2614
rect 2990 2610 3050 2614
rect 2990 1430 3050 1490
rect 655 1200 805 1350
rect 2995 1200 3145 1350
rect 3312 1122 3368 1178
<< metal3 >>
rect 1325 2690 1395 2695
rect 485 2670 555 2675
rect 485 2610 490 2670
rect 550 2610 555 2670
rect 1325 2630 1330 2690
rect 1390 2630 1395 2690
rect 1325 2625 1395 2630
rect 2095 2690 2165 2695
rect 2095 2630 2100 2690
rect 2160 2630 2165 2690
rect 2095 2625 2165 2630
rect 2985 2670 3055 2675
rect 485 2605 555 2610
rect 490 1130 550 2605
rect 650 1350 810 1355
rect 650 1345 655 1350
rect 805 1345 810 1350
rect 650 1189 810 1195
rect 420 850 550 1130
rect 1330 840 1390 2625
rect 2100 810 2160 2625
rect 2985 2610 2990 2670
rect 3050 2610 3055 2670
rect 2985 2605 3055 2610
rect 2990 1495 3050 2605
rect 2985 1490 3055 1495
rect 2985 1430 2990 1490
rect 3050 1430 3055 1490
rect 2985 1425 3055 1430
rect 2990 1350 3150 1355
rect 2990 1345 2995 1350
rect 3145 1345 3150 1350
rect 2990 1189 3150 1195
rect 3307 1178 3373 1183
rect 3307 1122 3312 1178
rect 3368 1122 3373 1178
rect 3307 1117 3373 1122
rect 3310 850 3370 1117
<< via3 >>
rect 650 1200 655 1345
rect 655 1200 805 1345
rect 805 1200 810 1345
rect 650 1195 810 1200
rect 2990 1200 2995 1345
rect 2995 1200 3145 1345
rect 3145 1200 3150 1345
rect 2990 1195 3150 1200
<< metal4 >>
rect 649 1345 811 1346
rect 649 1195 650 1345
rect 810 1195 811 1345
rect 649 1194 811 1195
rect 2989 1345 3151 1346
rect 2989 1195 2990 1345
rect 3150 1195 3151 1345
rect 2989 1194 3151 1195
rect 655 1115 805 1194
rect 660 410 740 1115
rect 2995 1055 3145 1194
rect 3050 430 3110 1055
rect 370 400 880 410
rect 280 340 960 400
rect 2650 370 3550 430
rect 370 330 880 340
use sky130_fd_pr__cap_mim_m3_1_9SN4GA  XC29
timestamp 1672355014
transform 0 -1 1265 1 0 411
box -610 -464 610 464
use sky130_fd_pr__cap_mim_m3_1_9SN4GA  XC30
timestamp 1672355014
transform 0 -1 2465 1 0 411
box -610 -464 610 464
use sky130_fd_pr__nfet_01v8_Q8AFGD  XM19
timestamp 1672367450
transform 1 0 -1187 0 1 1712
box -212 -310 212 310
use sky130_fd_pr__nfet_01v8_Q8AFGD  XM80
timestamp 1672367450
transform 1 0 -587 0 1 1712
box -212 -310 212 310
use sky130_fd_pr__pfet_01v8_8DZSMJ  XM81
timestamp 1672367450
transform 1 0 -587 0 1 4719
box -212 -319 212 319
use sky130_fd_pr__pfet_01v8_8DZSMJ  XM82
timestamp 1672367450
transform 1 0 232 0 1 4719
box -212 -319 212 319
use sky130_fd_pr__pfet_01v8_8DZSMJ  XM83
timestamp 1672367450
transform 1 0 213 0 1 3719
box -212 -319 212 319
use sky130_fd_pr__nfet_01v8_Q8AFGD  XM85
timestamp 1672367450
transform 1 0 213 0 1 1712
box -212 -310 212 310
use sky130_fd_pr__nfet_01v8_Q8AFGD  XM86
timestamp 1672367450
transform 1 0 213 0 1 2712
box -212 -310 212 310
use sky130_fd_pr__pfet_01v8_8DZSMJ  XM87
timestamp 1672367450
transform 1 0 1013 0 1 4719
box -212 -319 212 319
use sky130_fd_pr__pfet_01v8_8DZSMJ  XM88
timestamp 1672367450
transform 1 0 1013 0 1 3719
box -212 -319 212 319
use sky130_fd_pr__nfet_01v8_Q8AFGD  XM90
timestamp 1672367450
transform 1 0 1013 0 1 2712
box -212 -310 212 310
use sky130_fd_pr__nfet_01v8_Q8AFGD  XM91
timestamp 1672367450
transform 1 0 1013 0 1 1712
box -212 -310 212 310
use sky130_fd_pr__pfet_01v8_8DZSMJ  XM92
timestamp 1672367450
transform 1 0 1813 0 1 4719
box -212 -319 212 319
use sky130_fd_pr__pfet_01v8_8DZSMJ  XM93
timestamp 1672367450
transform 1 0 1813 0 1 3719
box -212 -319 212 319
use sky130_fd_pr__nfet_01v8_Q8AFGD  XM95
timestamp 1672367450
transform 1 0 1813 0 1 2712
box -212 -310 212 310
use sky130_fd_pr__nfet_01v8_Q8AFGD  XM96
timestamp 1672367450
transform 1 0 1813 0 1 1712
box -212 -310 212 310
use sky130_fd_pr__pfet_01v8_8DZSMJ  XM97
timestamp 1672367450
transform 1 0 2613 0 1 4719
box -212 -319 212 319
use sky130_fd_pr__pfet_01v8_8DZSMJ  XM98
timestamp 1672367450
transform 1 0 2613 0 1 3719
box -212 -319 212 319
use sky130_fd_pr__nfet_01v8_Q8AFGD  XM100
timestamp 1672367450
transform 1 0 2613 0 1 2712
box -212 -310 212 310
use sky130_fd_pr__pfet_01v8_8DZSMJ  XM102
timestamp 1672367450
transform 1 0 3413 0 1 4719
box -212 -319 212 319
use sky130_fd_pr__nfet_01v8_Q8AFGD  XM105
timestamp 1672367450
transform 1 0 3413 0 1 2712
box -212 -310 212 310
use sky130_fd_pr__pfet_01v8_lvt_D3C9B3  XM107
timestamp 1672367450
transform 1 0 -1967 0 1 5469
box -232 -269 232 269
use sky130_fd_pr__res_xhigh_po_0p69_ET3NLF  XR38
timestamp 1672367450
transform 1 0 -1965 0 1 3231
box -235 -1829 235 1829
use sky130_fd_pr__res_xhigh_po_0p35_H4KU7R  XR40
timestamp 1672367450
transform 1 0 -1199 0 1 4201
box -201 -1999 201 1999
use sky130_fd_pr__cap_mim_m3_1_9SN4GA  sky130_fd_pr__cap_mim_m3_1_9SN4GA_0
timestamp 1672355014
transform 0 -1 3665 1 0 411
box -610 -464 610 464
use sky130_fd_pr__cap_mim_m3_1_9SN4GA  sky130_fd_pr__cap_mim_m3_1_9SN4GA_1
timestamp 1672355014
transform 0 -1 65 1 0 411
box -610 -464 610 464
use sky130_fd_pr__nfet_01v8_Q8AFGD  sky130_fd_pr__nfet_01v8_Q8AFGD_0
timestamp 1672367450
transform 1 0 2613 0 1 1712
box -212 -310 212 310
use sky130_fd_pr__nfet_01v8_Q8AFGD  sky130_fd_pr__nfet_01v8_Q8AFGD_1
timestamp 1672367450
transform 1 0 3413 0 1 1712
box -212 -310 212 310
use sky130_fd_pr__pfet_01v8_8DZSMJ  sky130_fd_pr__pfet_01v8_8DZSMJ_0
timestamp 1672367450
transform 1 0 3413 0 1 3719
box -212 -319 212 319
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1669390400
transform -1 0 4716 0 -1 3600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  x4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1669390400
transform -1 0 4234 0 -1 3592
box -38 -48 314 592
<< labels >>
rlabel metal1 220 5160 290 5230 1 vcc
port 0 n
rlabel metal1 -1680 5330 -1650 5360 1 ctrl
port 1 n
rlabel metal1 1110 1240 1140 1270 1 gnd
port 2 n
rlabel locali 4308 3362 4320 3372 1 out
port 3 n
<< end >>
