magic
tech sky130A
magscale 1 2
timestamp 1672355014
<< metal3 >>
rect -612 437 612 465
rect -612 -437 528 437
rect 592 -437 612 437
rect -612 -465 612 -437
<< via3 >>
rect 528 -437 592 437
<< mimcap >>
rect -572 385 280 425
rect -572 -385 -532 385
rect 240 -385 280 385
rect -572 -425 280 -385
<< mimcapcontact >>
rect -532 -385 240 385
<< metal4 >>
rect 512 437 608 453
rect -533 385 241 386
rect -533 -385 -532 385
rect 240 -385 241 385
rect -533 -386 241 -385
rect 512 -437 528 437
rect 592 -437 608 437
rect 512 -453 608 -437
<< properties >>
string FIXED_BBOX -612 -465 320 465
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 4.255 l 4.25 val 39.399 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
