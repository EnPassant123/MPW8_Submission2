magic
tech sky130A
timestamp 1672028832
<< end >>
