magic
tech sky130A
magscale 1 2
timestamp 1672367450
<< error_p >>
rect -29 172 29 178
rect -29 138 -17 172
rect -29 132 29 138
rect -29 -138 29 -132
rect -29 -172 -17 -138
rect -29 -178 29 -172
<< pwell >>
rect -212 -310 212 310
<< nmos >>
rect -16 -100 16 100
<< ndiff >>
rect -74 88 -16 100
rect -74 -88 -62 88
rect -28 -88 -16 88
rect -74 -100 -16 -88
rect 16 88 74 100
rect 16 -88 28 88
rect 62 -88 74 88
rect 16 -100 74 -88
<< ndiffc >>
rect -62 -88 -28 88
rect 28 -88 62 88
<< psubdiff >>
rect -176 240 -80 274
rect 80 240 176 274
rect -176 178 -142 240
rect 142 178 176 240
rect -176 -240 -142 -178
rect 142 -240 176 -178
rect -176 -274 -80 -240
rect 80 -274 176 -240
<< psubdiffcont >>
rect -80 240 80 274
rect -176 -178 -142 178
rect 142 -178 176 178
rect -80 -274 80 -240
<< poly >>
rect -33 172 33 188
rect -33 138 -17 172
rect 17 138 33 172
rect -33 122 33 138
rect -16 100 16 122
rect -16 -122 16 -100
rect -33 -138 33 -122
rect -33 -172 -17 -138
rect 17 -172 33 -138
rect -33 -188 33 -172
<< polycont >>
rect -17 138 17 172
rect -17 -172 17 -138
<< locali >>
rect -176 240 -80 274
rect 80 240 176 274
rect -176 178 -142 240
rect 142 178 176 240
rect -33 138 -17 172
rect 17 138 33 172
rect -62 88 -28 104
rect -62 -104 -28 -88
rect 28 88 62 104
rect 28 -104 62 -88
rect -33 -172 -17 -138
rect 17 -172 33 -138
rect -176 -240 -142 -178
rect 142 -240 176 -178
rect -176 -274 -80 -240
rect 80 -274 176 -240
<< viali >>
rect -17 138 17 172
rect -62 -88 -28 88
rect 28 -88 62 88
rect -17 -172 17 -138
<< metal1 >>
rect -29 172 29 178
rect -29 138 -17 172
rect 17 138 29 172
rect -29 132 29 138
rect -68 88 -22 100
rect -68 -88 -62 88
rect -28 -88 -22 88
rect -68 -100 -22 -88
rect 22 88 68 100
rect 22 -88 28 88
rect 62 -88 68 88
rect 22 -100 68 -88
rect -29 -138 29 -132
rect -29 -172 -17 -138
rect 17 -172 29 -138
rect -29 -178 29 -172
<< properties >>
string FIXED_BBOX -159 -257 159 257
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 0.155 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
