magic
tech sky130A
timestamp 1671933972
<< pwell >>
rect -248 -1105 248 1105
<< nmos >>
rect -150 -1000 150 1000
<< ndiff >>
rect -179 994 -150 1000
rect -179 -994 -173 994
rect -156 -994 -150 994
rect -179 -1000 -150 -994
rect 150 994 179 1000
rect 150 -994 156 994
rect 173 -994 179 994
rect 150 -1000 179 -994
<< ndiffc >>
rect -173 -994 -156 994
rect 156 -994 173 994
<< psubdiff >>
rect -230 1070 -182 1087
rect 182 1070 230 1087
rect -230 1039 -213 1070
rect 213 1039 230 1070
rect -230 -1070 -213 -1039
rect 213 -1070 230 -1039
rect -230 -1087 -182 -1070
rect 182 -1087 230 -1070
<< psubdiffcont >>
rect -182 1070 182 1087
rect -230 -1039 -213 1039
rect 213 -1039 230 1039
rect -182 -1087 182 -1070
<< poly >>
rect -150 1036 150 1044
rect -150 1019 -142 1036
rect 142 1019 150 1036
rect -150 1000 150 1019
rect -150 -1019 150 -1000
rect -150 -1036 -142 -1019
rect 142 -1036 150 -1019
rect -150 -1044 150 -1036
<< polycont >>
rect -142 1019 142 1036
rect -142 -1036 142 -1019
<< locali >>
rect -230 1070 -182 1087
rect 182 1070 230 1087
rect -230 1039 -213 1070
rect 213 1039 230 1070
rect -150 1019 -142 1036
rect 142 1019 150 1036
rect -173 994 -156 1002
rect -173 -1002 -156 -994
rect 156 994 173 1002
rect 156 -1002 173 -994
rect -150 -1036 -142 -1019
rect 142 -1036 150 -1019
rect -230 -1070 -213 -1039
rect 213 -1070 230 -1039
rect -230 -1087 -182 -1070
rect 182 -1087 230 -1070
<< viali >>
rect -142 1019 142 1036
rect -173 -994 -156 994
rect 156 -994 173 994
rect -142 -1036 142 -1019
<< metal1 >>
rect -148 1036 148 1039
rect -148 1019 -142 1036
rect 142 1019 148 1036
rect -148 1016 148 1019
rect -176 994 -153 1000
rect -176 -994 -173 994
rect -156 -994 -153 994
rect -176 -1000 -153 -994
rect 153 994 176 1000
rect 153 -994 156 994
rect 173 -994 176 994
rect 153 -1000 176 -994
rect -148 -1019 148 -1016
rect -148 -1036 -142 -1019
rect 142 -1036 148 -1019
rect -148 -1039 148 -1036
<< properties >>
string FIXED_BBOX -221 -1078 221 1078
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 20 l 3 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
