magic
tech sky130A
magscale 1 2
timestamp 1672362834
<< pwell >>
rect -247 -1210 247 1210
<< nmos >>
rect -51 -1000 51 1000
<< ndiff >>
rect -109 988 -51 1000
rect -109 -988 -97 988
rect -63 -988 -51 988
rect -109 -1000 -51 -988
rect 51 988 109 1000
rect 51 -988 63 988
rect 97 -988 109 988
rect 51 -1000 109 -988
<< ndiffc >>
rect -97 -988 -63 988
rect 63 -988 97 988
<< psubdiff >>
rect -211 1140 -115 1174
rect 115 1140 211 1174
rect -211 1078 -177 1140
rect 177 1078 211 1140
rect -211 -1140 -177 -1078
rect 177 -1140 211 -1078
rect -211 -1174 -115 -1140
rect 115 -1174 211 -1140
<< psubdiffcont >>
rect -115 1140 115 1174
rect -211 -1078 -177 1078
rect 177 -1078 211 1078
rect -115 -1174 115 -1140
<< poly >>
rect -51 1072 51 1088
rect -51 1038 -35 1072
rect 35 1038 51 1072
rect -51 1000 51 1038
rect -51 -1038 51 -1000
rect -51 -1072 -35 -1038
rect 35 -1072 51 -1038
rect -51 -1088 51 -1072
<< polycont >>
rect -35 1038 35 1072
rect -35 -1072 35 -1038
<< locali >>
rect -211 1140 -115 1174
rect 115 1140 211 1174
rect -211 1078 -177 1140
rect 177 1078 211 1140
rect -51 1038 -35 1072
rect 35 1038 51 1072
rect -97 988 -63 1004
rect -97 -1004 -63 -988
rect 63 988 97 1004
rect 63 -1004 97 -988
rect -51 -1072 -35 -1038
rect 35 -1072 51 -1038
rect -211 -1140 -177 -1078
rect 177 -1140 211 -1078
rect -211 -1174 -115 -1140
rect 115 -1174 211 -1140
<< viali >>
rect -35 1038 35 1072
rect -97 -988 -63 988
rect 63 -988 97 988
rect -35 -1072 35 -1038
<< metal1 >>
rect -47 1072 47 1078
rect -47 1038 -35 1072
rect 35 1038 47 1072
rect -47 1032 47 1038
rect -103 988 -57 1000
rect -103 -988 -97 988
rect -63 -988 -57 988
rect -103 -1000 -57 -988
rect 57 988 103 1000
rect 57 -988 63 988
rect 97 -988 103 988
rect 57 -1000 103 -988
rect -47 -1038 47 -1032
rect -47 -1072 -35 -1038
rect 35 -1072 47 -1038
rect -47 -1078 47 -1072
<< properties >>
string FIXED_BBOX -194 -1157 194 1157
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 10 l 0.505 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
