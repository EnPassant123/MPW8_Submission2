magic
tech sky130A
timestamp 1672007445
<< pwell >>
rect -100 -1799 100 1799
<< psubdiff >>
rect -82 1764 -34 1781
rect 34 1764 82 1781
rect -82 1733 -65 1764
rect 65 1733 82 1764
rect -82 -1764 -65 -1733
rect 65 -1764 82 -1733
rect -82 -1781 -34 -1764
rect 34 -1781 82 -1764
<< psubdiffcont >>
rect -34 1764 34 1781
rect -82 -1733 -65 1733
rect 65 -1733 82 1733
rect -34 -1781 34 -1764
<< xpolycontact >>
rect -17 1500 17 1716
rect -17 -1716 17 -1500
<< xpolyres >>
rect -17 -1500 17 1500
<< locali >>
rect -82 1764 -34 1781
rect 34 1764 82 1781
rect -82 1733 -65 1764
rect 65 1733 82 1764
rect -82 -1764 -65 -1733
rect 65 -1764 82 -1733
rect -82 -1781 -34 -1764
rect 34 -1781 82 -1764
<< viali >>
rect -9 1508 9 1707
rect -9 -1707 9 -1508
<< metal1 >>
rect -12 1707 12 1713
rect -12 1508 -9 1707
rect 9 1508 12 1707
rect -12 1502 12 1508
rect -12 -1508 12 -1502
rect -12 -1707 -9 -1508
rect 9 -1707 12 -1508
rect -12 -1713 12 -1707
<< res0p35 >>
rect -18 -1501 18 1501
<< properties >>
string FIXED_BBOX -74 -1772 74 1772
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 30 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 172.504k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
