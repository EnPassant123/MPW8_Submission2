magic
tech sky130A
magscale 1 2
timestamp 1672468335
<< pwell >>
rect -497 -2210 497 2210
<< nmos >>
rect -301 -2000 301 2000
<< ndiff >>
rect -359 1988 -301 2000
rect -359 -1988 -347 1988
rect -313 -1988 -301 1988
rect -359 -2000 -301 -1988
rect 301 1988 359 2000
rect 301 -1988 313 1988
rect 347 -1988 359 1988
rect 301 -2000 359 -1988
<< ndiffc >>
rect -347 -1988 -313 1988
rect 313 -1988 347 1988
<< psubdiff >>
rect -461 2140 -365 2174
rect 365 2140 461 2174
rect -461 2078 -427 2140
rect 427 2078 461 2140
rect -461 -2140 -427 -2078
rect 427 -2140 461 -2078
rect -461 -2174 -365 -2140
rect 365 -2174 461 -2140
<< psubdiffcont >>
rect -365 2140 365 2174
rect -461 -2078 -427 2078
rect 427 -2078 461 2078
rect -365 -2174 365 -2140
<< poly >>
rect -301 2072 301 2088
rect -301 2038 -285 2072
rect 285 2038 301 2072
rect -301 2000 301 2038
rect -301 -2038 301 -2000
rect -301 -2072 -285 -2038
rect 285 -2072 301 -2038
rect -301 -2088 301 -2072
<< polycont >>
rect -285 2038 285 2072
rect -285 -2072 285 -2038
<< locali >>
rect -461 2140 -365 2174
rect 365 2140 461 2174
rect -461 2078 -427 2140
rect 427 2078 461 2140
rect -301 2038 -285 2072
rect 285 2038 301 2072
rect -347 1988 -313 2004
rect -347 -2004 -313 -1988
rect 313 1988 347 2004
rect 313 -2004 347 -1988
rect -301 -2072 -285 -2038
rect 285 -2072 301 -2038
rect -461 -2140 -427 -2078
rect 427 -2140 461 -2078
rect -461 -2174 -365 -2140
rect 365 -2174 461 -2140
<< viali >>
rect -285 2038 285 2072
rect -347 -1988 -313 1988
rect 313 -1988 347 1988
rect -285 -2072 285 -2038
<< metal1 >>
rect -297 2072 297 2078
rect -297 2038 -285 2072
rect 285 2038 297 2072
rect -297 2032 297 2038
rect -353 1988 -307 2000
rect -353 -1988 -347 1988
rect -313 -1988 -307 1988
rect -353 -2000 -307 -1988
rect 307 1988 353 2000
rect 307 -1988 313 1988
rect 347 -1988 353 1988
rect 307 -2000 353 -1988
rect -297 -2038 297 -2032
rect -297 -2072 -285 -2038
rect 285 -2072 297 -2038
rect -297 -2078 297 -2072
<< properties >>
string FIXED_BBOX -444 -2157 444 2157
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 20 l 3.005 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
