magic
tech sky130A
timestamp 1672354625
<< pwell >>
rect -123 -3055 123 3055
<< nmoslvt >>
rect -25 -2950 25 2950
<< ndiff >>
rect -54 2944 -25 2950
rect -54 -2944 -48 2944
rect -31 -2944 -25 2944
rect -54 -2950 -25 -2944
rect 25 2944 54 2950
rect 25 -2944 31 2944
rect 48 -2944 54 2944
rect 25 -2950 54 -2944
<< ndiffc >>
rect -48 -2944 -31 2944
rect 31 -2944 48 2944
<< psubdiff >>
rect -105 3020 -57 3037
rect 57 3020 105 3037
rect -105 2989 -88 3020
rect 88 2989 105 3020
rect -105 -3020 -88 -2989
rect 88 -3020 105 -2989
rect -105 -3037 -57 -3020
rect 57 -3037 105 -3020
<< psubdiffcont >>
rect -57 3020 57 3037
rect -105 -2989 -88 2989
rect 88 -2989 105 2989
rect -57 -3037 57 -3020
<< poly >>
rect -25 2986 25 2994
rect -25 2969 -17 2986
rect 17 2969 25 2986
rect -25 2950 25 2969
rect -25 -2969 25 -2950
rect -25 -2986 -17 -2969
rect 17 -2986 25 -2969
rect -25 -2994 25 -2986
<< polycont >>
rect -17 2969 17 2986
rect -17 -2986 17 -2969
<< locali >>
rect -105 3020 -57 3037
rect 57 3020 105 3037
rect -105 2989 -88 3020
rect 88 2989 105 3020
rect -25 2969 -17 2986
rect 17 2969 25 2986
rect -48 2944 -31 2952
rect -48 -2952 -31 -2944
rect 31 2944 48 2952
rect 31 -2952 48 -2944
rect -25 -2986 -17 -2969
rect 17 -2986 25 -2969
rect -105 -3020 -88 -2989
rect 88 -3020 105 -2989
rect -105 -3037 -57 -3020
rect 57 -3037 105 -3020
<< viali >>
rect -17 2969 17 2986
rect -48 -2944 -31 2944
rect 31 -2944 48 2944
rect -17 -2986 17 -2969
<< metal1 >>
rect -23 2986 23 2989
rect -23 2969 -17 2986
rect 17 2969 23 2986
rect -23 2966 23 2969
rect -51 2944 -28 2950
rect -51 -2944 -48 2944
rect -31 -2944 -28 2944
rect -51 -2950 -28 -2944
rect 28 2944 51 2950
rect 28 -2944 31 2944
rect 48 -2944 51 2944
rect 28 -2950 51 -2944
rect -23 -2969 23 -2966
rect -23 -2986 -17 -2969
rect 17 -2986 23 -2969
rect -23 -2989 23 -2986
<< properties >>
string FIXED_BBOX -96 -3028 96 3028
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 59.0 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
