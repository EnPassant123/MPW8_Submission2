magic
tech sky130A
magscale 1 2
timestamp 1672370185
<< pwell >>
rect -201 -1469 201 1469
<< psubdiff >>
rect -165 1399 -69 1433
rect 69 1399 165 1433
rect -165 1337 -131 1399
rect 131 1337 165 1399
rect -165 -1399 -131 -1337
rect 131 -1399 165 -1337
rect -165 -1433 -69 -1399
rect 69 -1433 165 -1399
<< psubdiffcont >>
rect -69 1399 69 1433
rect -165 -1337 -131 1337
rect 131 -1337 165 1337
rect -69 -1433 69 -1399
<< xpolycontact >>
rect -35 871 35 1303
rect -35 -1303 35 -871
<< xpolyres >>
rect -35 -871 35 871
<< locali >>
rect -165 1399 -69 1433
rect 69 1399 165 1433
rect -165 1337 -131 1399
rect 131 1337 165 1399
rect -165 -1399 -131 -1337
rect 131 -1399 165 -1337
rect -165 -1433 -69 -1399
rect 69 -1433 165 -1399
<< viali >>
rect -19 888 19 1285
rect -19 -1285 19 -888
<< metal1 >>
rect -25 1285 25 1297
rect -25 888 -19 1285
rect 19 888 25 1285
rect -25 876 25 888
rect -25 -888 25 -876
rect -25 -1285 -19 -888
rect 19 -1285 25 -888
rect -25 -1297 25 -1285
<< res0p35 >>
rect -37 -873 37 873
<< properties >>
string FIXED_BBOX -148 -1416 148 1416
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 8.705 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 50.818k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
