magic
tech sky130A
magscale 1 2
timestamp 1672368307
<< nwell >>
rect -247 -1219 247 1219
<< pmos >>
rect -51 -1000 51 1000
<< pdiff >>
rect -109 988 -51 1000
rect -109 -988 -97 988
rect -63 -988 -51 988
rect -109 -1000 -51 -988
rect 51 988 109 1000
rect 51 -988 63 988
rect 97 -988 109 988
rect 51 -1000 109 -988
<< pdiffc >>
rect -97 -988 -63 988
rect 63 -988 97 988
<< nsubdiff >>
rect -211 1149 -115 1183
rect 115 1149 211 1183
rect -211 1087 -177 1149
rect 177 1087 211 1149
rect -211 -1149 -177 -1087
rect 177 -1149 211 -1087
rect -211 -1183 -115 -1149
rect 115 -1183 211 -1149
<< nsubdiffcont >>
rect -115 1149 115 1183
rect -211 -1087 -177 1087
rect 177 -1087 211 1087
rect -115 -1183 115 -1149
<< poly >>
rect -51 1081 51 1097
rect -51 1047 -35 1081
rect 35 1047 51 1081
rect -51 1000 51 1047
rect -51 -1047 51 -1000
rect -51 -1081 -35 -1047
rect 35 -1081 51 -1047
rect -51 -1097 51 -1081
<< polycont >>
rect -35 1047 35 1081
rect -35 -1081 35 -1047
<< locali >>
rect -211 1149 -115 1183
rect 115 1149 211 1183
rect -211 1087 -177 1149
rect 177 1087 211 1149
rect -51 1047 -35 1081
rect 35 1047 51 1081
rect -97 988 -63 1004
rect -97 -1004 -63 -988
rect 63 988 97 1004
rect 63 -1004 97 -988
rect -51 -1081 -35 -1047
rect 35 -1081 51 -1047
rect -211 -1149 -177 -1087
rect 177 -1149 211 -1087
rect -211 -1183 -115 -1149
rect 115 -1183 211 -1149
<< viali >>
rect -35 1047 35 1081
rect -97 -988 -63 988
rect 63 -988 97 988
rect -35 -1081 35 -1047
<< metal1 >>
rect -47 1081 47 1087
rect -47 1047 -35 1081
rect 35 1047 47 1081
rect -47 1041 47 1047
rect -103 988 -57 1000
rect -103 -988 -97 988
rect -63 -988 -57 988
rect -103 -1000 -57 -988
rect 57 988 103 1000
rect 57 -988 63 988
rect 97 -988 103 988
rect 57 -1000 103 -988
rect -47 -1047 47 -1041
rect -47 -1081 -35 -1047
rect 35 -1081 47 -1047
rect -47 -1087 47 -1081
<< properties >>
string FIXED_BBOX -194 -1166 194 1166
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 10 l 0.505 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
